*** Fig 2. Circuitfile 

.model jj0 jj(rtype=0, icrit=5.0000uA, cap=60.0000fF) 
*SQUID embedded transmission line 
Ip 0 1 sin(0 5.7000uA 12.0000GHz 9ns 0 0)
Is 0 1 sin(0 0.3000uA 7.2000GHz 9ns 0 0) 

Vmeas0 1 2 0V
Rtermfront 2 0 23.8747Ohm
Vmeas1 2 3 0V

*Flux Biasing 
Idc2 0 50002 pwl(0 0uA 5ns 14.0680uA) 
Lflux2 50002 0 57.0000pH 
K2 Lg2 Lflux2 1

Cg2 3 0 50.0000fF 
Lg2 3 4 57.0000pH
B2 3 4 10001 jj0 
Cgg2 4 0 50.0000fF
Vmeas2 4 5 0V

*Flux Biasing 
Idc3 0 50003 pwl(0 0uA 5ns 14.0680uA) 
Lflux3 50003 0 57.0000pH 
K3 Lg3 Lflux3 1

Cg3 5 0 50.0000fF 
Lg3 5 6 57.0000pH
B3 5 6 10002 jj0 
Cgg3 6 0 50.0000fF
Vmeas3 6 7 0V

*Flux Biasing 
Idc4 0 50004 pwl(0 0uA 5ns 14.0680uA) 
Lflux4 50004 0 57.0000pH 
K4 Lg4 Lflux4 1

Cg4 7 0 50.0000fF 
Lg4 7 8 57.0000pH
B4 7 8 10003 jj0 
Cgg4 8 0 50.0000fF
Vmeas4 8 9 0V

*Flux Biasing 
Idc5 0 50005 pwl(0 0uA 5ns 14.0680uA) 
Lflux5 50005 0 57.0000pH 
K5 Lg5 Lflux5 1

Cg5 9 0 50.0000fF 
Lg5 9 10 57.0000pH
B5 9 10 10004 jj0 
Cgg5 10 0 50.0000fF
Vmeas5 10 11 0V

*Flux Biasing 
Idc6 0 50006 pwl(0 0uA 5ns 14.0680uA) 
Lflux6 50006 0 57.0000pH 
K6 Lg6 Lflux6 1

Cg6 11 0 50.0000fF 
Lg6 11 12 57.0000pH
B6 11 12 10005 jj0 
Cgg6 12 0 50.0000fF
Vmeas6 12 13 0V

*Flux Biasing 
Idc7 0 50007 pwl(0 0uA 5ns 14.0680uA) 
Lflux7 50007 0 57.0000pH 
K7 Lg7 Lflux7 1

Cg7 13 0 50.0000fF 
Lg7 13 14 57.0000pH
B7 13 14 10006 jj0 
Cgg7 14 0 50.0000fF
Vmeas7 14 15 0V

*Flux Biasing 
Idc8 0 50008 pwl(0 0uA 5ns 14.0680uA) 
Lflux8 50008 0 57.0000pH 
K8 Lg8 Lflux8 1

Cg8 15 0 50.0000fF 
Lg8 15 16 57.0000pH
B8 15 16 10007 jj0 
Cgg8 16 0 50.0000fF
Vmeas8 16 17 0V

*Flux Biasing 
Idc9 0 50009 pwl(0 0uA 5ns 14.0680uA) 
Lflux9 50009 0 57.0000pH 
K9 Lg9 Lflux9 1

Cg9 17 0 50.0000fF 
Lg9 17 18 57.0000pH
B9 17 18 10008 jj0 
Cgg9 18 0 50.0000fF
Vmeas9 18 19 0V

*Flux Biasing 
Idc10 0 50010 pwl(0 0uA 5ns 14.0680uA) 
Lflux10 50010 0 57.0000pH 
K10 Lg10 Lflux10 1

Cg10 19 0 50.0000fF 
Lg10 19 20 57.0000pH
B10 19 20 10009 jj0 
Cgg10 20 0 50.0000fF
Vmeas10 20 21 0V

*Flux Biasing 
Idc11 0 50011 pwl(0 0uA 5ns 14.0680uA) 
Lflux11 50011 0 57.0000pH 
K11 Lg11 Lflux11 1

Cg11 21 0 50.0000fF 
Lg11 21 22 57.0000pH
B11 21 22 10010 jj0 
Cgg11 22 0 50.0000fF
Vmeas11 22 23 0V

*Flux Biasing 
Idc12 0 50012 pwl(0 0uA 5ns 14.0680uA) 
Lflux12 50012 0 57.0000pH 
K12 Lg12 Lflux12 1

Cg12 23 0 50.0000fF 
Lg12 23 24 57.0000pH
B12 23 24 10011 jj0 
Cgg12 24 0 50.0000fF
Vmeas12 24 25 0V

*Flux Biasing 
Idc13 0 50013 pwl(0 0uA 5ns 14.0680uA) 
Lflux13 50013 0 57.0000pH 
K13 Lg13 Lflux13 1

Cg13 25 0 50.0000fF 
Lg13 25 26 57.0000pH
B13 25 26 10012 jj0 
Cgg13 26 0 50.0000fF
Vmeas13 26 27 0V

*Flux Biasing 
Idc14 0 50014 pwl(0 0uA 5ns 14.0680uA) 
Lflux14 50014 0 57.0000pH 
K14 Lg14 Lflux14 1

Cg14 27 0 50.0000fF 
Lg14 27 28 57.0000pH
B14 27 28 10013 jj0 
Cgg14 28 0 50.0000fF
Vmeas14 28 29 0V

*Flux Biasing 
Idc15 0 50015 pwl(0 0uA 5ns 14.0680uA) 
Lflux15 50015 0 57.0000pH 
K15 Lg15 Lflux15 1

Cg15 29 0 50.0000fF 
Lg15 29 30 57.0000pH
B15 29 30 10014 jj0 
Cgg15 30 0 50.0000fF
Vmeas15 30 31 0V

*Flux Biasing 
Idc16 0 50016 pwl(0 0uA 5ns 14.0680uA) 
Lflux16 50016 0 57.0000pH 
K16 Lg16 Lflux16 1

Cg16 31 0 50.0000fF 
Lg16 31 32 57.0000pH
B16 31 32 10015 jj0 
Cgg16 32 0 50.0000fF
Vmeas16 32 33 0V

*Flux Biasing 
Idc17 0 50017 pwl(0 0uA 5ns 14.0680uA) 
Lflux17 50017 0 57.0000pH 
K17 Lg17 Lflux17 1

Cg17 33 0 50.0000fF 
Lg17 33 34 57.0000pH
B17 33 34 10016 jj0 
Cgg17 34 0 50.0000fF
Vmeas17 34 35 0V

*Flux Biasing 
Idc18 0 50018 pwl(0 0uA 5ns 14.0680uA) 
Lflux18 50018 0 57.0000pH 
K18 Lg18 Lflux18 1

Cg18 35 0 50.0000fF 
Lg18 35 36 57.0000pH
B18 35 36 10017 jj0 
Cgg18 36 0 50.0000fF
Vmeas18 36 37 0V

*Flux Biasing 
Idc19 0 50019 pwl(0 0uA 5ns 14.0680uA) 
Lflux19 50019 0 57.0000pH 
K19 Lg19 Lflux19 1

Cg19 37 0 50.0000fF 
Lg19 37 38 57.0000pH
B19 37 38 10018 jj0 
Cgg19 38 0 50.0000fF
Vmeas19 38 39 0V

*Flux Biasing 
Idc20 0 50020 pwl(0 0uA 5ns 14.0680uA) 
Lflux20 50020 0 57.0000pH 
K20 Lg20 Lflux20 1

Cg20 39 0 50.0000fF 
Lg20 39 40 57.0000pH
B20 39 40 10019 jj0 
Cgg20 40 0 50.0000fF
Vmeas20 40 41 0V

*Flux Biasing 
Idc21 0 50021 pwl(0 0uA 5ns 14.0680uA) 
Lflux21 50021 0 57.0000pH 
K21 Lg21 Lflux21 1

Cg21 41 0 50.0000fF 
Lg21 41 42 57.0000pH
B21 41 42 10020 jj0 
Cgg21 42 0 50.0000fF
Vmeas21 42 43 0V

*Flux Biasing 
Idc22 0 50022 pwl(0 0uA 5ns 14.0680uA) 
Lflux22 50022 0 57.0000pH 
K22 Lg22 Lflux22 1

Cg22 43 0 50.0000fF 
Lg22 43 44 57.0000pH
B22 43 44 10021 jj0 
Cgg22 44 0 50.0000fF
Vmeas22 44 45 0V

*Flux Biasing 
Idc23 0 50023 pwl(0 0uA 5ns 14.0680uA) 
Lflux23 50023 0 57.0000pH 
K23 Lg23 Lflux23 1

Cg23 45 0 50.0000fF 
Lg23 45 46 57.0000pH
B23 45 46 10022 jj0 
Cgg23 46 0 50.0000fF
Vmeas23 46 47 0V

*Flux Biasing 
Idc24 0 50024 pwl(0 0uA 5ns 14.0680uA) 
Lflux24 50024 0 57.0000pH 
K24 Lg24 Lflux24 1

Cg24 47 0 50.0000fF 
Lg24 47 48 57.0000pH
B24 47 48 10023 jj0 
Cgg24 48 0 50.0000fF
Vmeas24 48 49 0V

*Flux Biasing 
Idc25 0 50025 pwl(0 0uA 5ns 14.0680uA) 
Lflux25 50025 0 57.0000pH 
K25 Lg25 Lflux25 1

Cg25 49 0 50.0000fF 
Lg25 49 50 57.0000pH
B25 49 50 10024 jj0 
Cgg25 50 0 50.0000fF
Vmeas25 50 51 0V

*Flux Biasing 
Idc26 0 50026 pwl(0 0uA 5ns 14.0680uA) 
Lflux26 50026 0 57.0000pH 
K26 Lg26 Lflux26 1

Cg26 51 0 50.0000fF 
Lg26 51 52 57.0000pH
B26 51 52 10025 jj0 
Cgg26 52 0 50.0000fF
Vmeas26 52 53 0V

*Flux Biasing 
Idc27 0 50027 pwl(0 0uA 5ns 14.0680uA) 
Lflux27 50027 0 57.0000pH 
K27 Lg27 Lflux27 1

Cg27 53 0 50.0000fF 
Lg27 53 54 57.0000pH
B27 53 54 10026 jj0 
Cgg27 54 0 50.0000fF
Vmeas27 54 55 0V

*Flux Biasing 
Idc28 0 50028 pwl(0 0uA 5ns 14.0680uA) 
Lflux28 50028 0 57.0000pH 
K28 Lg28 Lflux28 1

Cg28 55 0 50.0000fF 
Lg28 55 56 57.0000pH
B28 55 56 10027 jj0 
Cgg28 56 0 50.0000fF
Vmeas28 56 57 0V

*Flux Biasing 
Idc29 0 50029 pwl(0 0uA 5ns 14.0680uA) 
Lflux29 50029 0 57.0000pH 
K29 Lg29 Lflux29 1

Cg29 57 0 50.0000fF 
Lg29 57 58 57.0000pH
B29 57 58 10028 jj0 
Cgg29 58 0 50.0000fF
Vmeas29 58 59 0V

*Flux Biasing 
Idc30 0 50030 pwl(0 0uA 5ns 14.0680uA) 
Lflux30 50030 0 57.0000pH 
K30 Lg30 Lflux30 1

Cg30 59 0 50.0000fF 
Lg30 59 60 57.0000pH
B30 59 60 10029 jj0 
Cgg30 60 0 50.0000fF
Vmeas30 60 61 0V

*Flux Biasing 
Idc31 0 50031 pwl(0 0uA 5ns 14.0680uA) 
Lflux31 50031 0 57.0000pH 
K31 Lg31 Lflux31 1

Cg31 61 0 50.0000fF 
Lg31 61 62 57.0000pH
B31 61 62 10030 jj0 
Cgg31 62 0 50.0000fF
Vmeas31 62 63 0V

*Flux Biasing 
Idc32 0 50032 pwl(0 0uA 5ns 14.0680uA) 
Lflux32 50032 0 57.0000pH 
K32 Lg32 Lflux32 1

Cg32 63 0 50.0000fF 
Lg32 63 64 57.0000pH
B32 63 64 10031 jj0 
Cgg32 64 0 50.0000fF
Vmeas32 64 65 0V

*Flux Biasing 
Idc33 0 50033 pwl(0 0uA 5ns 14.0680uA) 
Lflux33 50033 0 57.0000pH 
K33 Lg33 Lflux33 1

Cg33 65 0 50.0000fF 
Lg33 65 66 57.0000pH
B33 65 66 10032 jj0 
Cgg33 66 0 50.0000fF
Vmeas33 66 67 0V

*Flux Biasing 
Idc34 0 50034 pwl(0 0uA 5ns 14.0680uA) 
Lflux34 50034 0 57.0000pH 
K34 Lg34 Lflux34 1

Cg34 67 0 50.0000fF 
Lg34 67 68 57.0000pH
B34 67 68 10033 jj0 
Cgg34 68 0 50.0000fF
Vmeas34 68 69 0V

*Flux Biasing 
Idc35 0 50035 pwl(0 0uA 5ns 14.0680uA) 
Lflux35 50035 0 57.0000pH 
K35 Lg35 Lflux35 1

Cg35 69 0 50.0000fF 
Lg35 69 70 57.0000pH
B35 69 70 10034 jj0 
Cgg35 70 0 50.0000fF
Vmeas35 70 71 0V

*Flux Biasing 
Idc36 0 50036 pwl(0 0uA 5ns 14.0680uA) 
Lflux36 50036 0 57.0000pH 
K36 Lg36 Lflux36 1

Cg36 71 0 50.0000fF 
Lg36 71 72 57.0000pH
B36 71 72 10035 jj0 
Cgg36 72 0 50.0000fF
Vmeas36 72 73 0V

*Flux Biasing 
Idc37 0 50037 pwl(0 0uA 5ns 14.0680uA) 
Lflux37 50037 0 57.0000pH 
K37 Lg37 Lflux37 1

Cg37 73 0 50.0000fF 
Lg37 73 74 57.0000pH
B37 73 74 10036 jj0 
Cgg37 74 0 50.0000fF
Vmeas37 74 75 0V

*Flux Biasing 
Idc38 0 50038 pwl(0 0uA 5ns 14.0680uA) 
Lflux38 50038 0 57.0000pH 
K38 Lg38 Lflux38 1

Cg38 75 0 50.0000fF 
Lg38 75 76 57.0000pH
B38 75 76 10037 jj0 
Cgg38 76 0 50.0000fF
Vmeas38 76 77 0V

*Flux Biasing 
Idc39 0 50039 pwl(0 0uA 5ns 14.0680uA) 
Lflux39 50039 0 57.0000pH 
K39 Lg39 Lflux39 1

Cg39 77 0 50.0000fF 
Lg39 77 78 57.0000pH
B39 77 78 10038 jj0 
Cgg39 78 0 50.0000fF
Vmeas39 78 79 0V

*Flux Biasing 
Idc40 0 50040 pwl(0 0uA 5ns 14.0680uA) 
Lflux40 50040 0 57.0000pH 
K40 Lg40 Lflux40 1

Cg40 79 0 50.0000fF 
Lg40 79 80 57.0000pH
B40 79 80 10039 jj0 
Cgg40 80 0 50.0000fF
Vmeas40 80 81 0V

*Flux Biasing 
Idc41 0 50041 pwl(0 0uA 5ns 14.0680uA) 
Lflux41 50041 0 57.0000pH 
K41 Lg41 Lflux41 1

Cg41 81 0 50.0000fF 
Lg41 81 82 57.0000pH
B41 81 82 10040 jj0 
Cgg41 82 0 50.0000fF
Vmeas41 82 83 0V

*Flux Biasing 
Idc42 0 50042 pwl(0 0uA 5ns 14.0680uA) 
Lflux42 50042 0 57.0000pH 
K42 Lg42 Lflux42 1

Cg42 83 0 50.0000fF 
Lg42 83 84 57.0000pH
B42 83 84 10041 jj0 
Cgg42 84 0 50.0000fF
Vmeas42 84 85 0V

*Flux Biasing 
Idc43 0 50043 pwl(0 0uA 5ns 14.0680uA) 
Lflux43 50043 0 57.0000pH 
K43 Lg43 Lflux43 1

Cg43 85 0 50.0000fF 
Lg43 85 86 57.0000pH
B43 85 86 10042 jj0 
Cgg43 86 0 50.0000fF
Vmeas43 86 87 0V

*Flux Biasing 
Idc44 0 50044 pwl(0 0uA 5ns 14.0680uA) 
Lflux44 50044 0 57.0000pH 
K44 Lg44 Lflux44 1

Cg44 87 0 50.0000fF 
Lg44 87 88 57.0000pH
B44 87 88 10043 jj0 
Cgg44 88 0 50.0000fF
Vmeas44 88 89 0V

*Flux Biasing 
Idc45 0 50045 pwl(0 0uA 5ns 14.0680uA) 
Lflux45 50045 0 57.0000pH 
K45 Lg45 Lflux45 1

Cg45 89 0 50.0000fF 
Lg45 89 90 57.0000pH
B45 89 90 10044 jj0 
Cgg45 90 0 50.0000fF
Vmeas45 90 91 0V

*Flux Biasing 
Idc46 0 50046 pwl(0 0uA 5ns 14.0680uA) 
Lflux46 50046 0 57.0000pH 
K46 Lg46 Lflux46 1

Cg46 91 0 50.0000fF 
Lg46 91 92 57.0000pH
B46 91 92 10045 jj0 
Cgg46 92 0 50.0000fF
Vmeas46 92 93 0V

*Flux Biasing 
Idc47 0 50047 pwl(0 0uA 5ns 14.0680uA) 
Lflux47 50047 0 57.0000pH 
K47 Lg47 Lflux47 1

Cg47 93 0 50.0000fF 
Lg47 93 94 57.0000pH
B47 93 94 10046 jj0 
Cgg47 94 0 50.0000fF
Vmeas47 94 95 0V

*Flux Biasing 
Idc48 0 50048 pwl(0 0uA 5ns 14.0680uA) 
Lflux48 50048 0 57.0000pH 
K48 Lg48 Lflux48 1

Cg48 95 0 50.0000fF 
Lg48 95 96 57.0000pH
B48 95 96 10047 jj0 
Cgg48 96 0 50.0000fF
Vmeas48 96 97 0V

*Flux Biasing 
Idc49 0 50049 pwl(0 0uA 5ns 14.0680uA) 
Lflux49 50049 0 57.0000pH 
K49 Lg49 Lflux49 1

Cg49 97 0 50.0000fF 
Lg49 97 98 57.0000pH
B49 97 98 10048 jj0 
Cgg49 98 0 50.0000fF
Vmeas49 98 99 0V

*Flux Biasing 
Idc50 0 50050 pwl(0 0uA 5ns 14.0680uA) 
Lflux50 50050 0 57.0000pH 
K50 Lg50 Lflux50 1

Cg50 99 0 50.0000fF 
Lg50 99 100 57.0000pH
B50 99 100 10049 jj0 
Cgg50 100 0 50.0000fF
Vmeas50 100 101 0V

*Flux Biasing 
Idc51 0 50051 pwl(0 0uA 5ns 14.0680uA) 
Lflux51 50051 0 57.0000pH 
K51 Lg51 Lflux51 1

Cg51 101 0 50.0000fF 
Lg51 101 102 57.0000pH
B51 101 102 10050 jj0 
Cgg51 102 0 50.0000fF
Vmeas51 102 103 0V

*Flux Biasing 
Idc52 0 50052 pwl(0 0uA 5ns 14.0680uA) 
Lflux52 50052 0 57.0000pH 
K52 Lg52 Lflux52 1

Cg52 103 0 50.0000fF 
Lg52 103 104 57.0000pH
B52 103 104 10051 jj0 
Cgg52 104 0 50.0000fF
Vmeas52 104 105 0V

*Flux Biasing 
Idc53 0 50053 pwl(0 0uA 5ns 14.0680uA) 
Lflux53 50053 0 57.0000pH 
K53 Lg53 Lflux53 1

Cg53 105 0 50.0000fF 
Lg53 105 106 57.0000pH
B53 105 106 10052 jj0 
Cgg53 106 0 50.0000fF
Vmeas53 106 107 0V

*Flux Biasing 
Idc54 0 50054 pwl(0 0uA 5ns 14.0680uA) 
Lflux54 50054 0 57.0000pH 
K54 Lg54 Lflux54 1

Cg54 107 0 50.0000fF 
Lg54 107 108 57.0000pH
B54 107 108 10053 jj0 
Cgg54 108 0 50.0000fF
Vmeas54 108 109 0V

*Flux Biasing 
Idc55 0 50055 pwl(0 0uA 5ns 14.0680uA) 
Lflux55 50055 0 57.0000pH 
K55 Lg55 Lflux55 1

Cg55 109 0 50.0000fF 
Lg55 109 110 57.0000pH
B55 109 110 10054 jj0 
Cgg55 110 0 50.0000fF
Vmeas55 110 111 0V

*Flux Biasing 
Idc56 0 50056 pwl(0 0uA 5ns 14.0680uA) 
Lflux56 50056 0 57.0000pH 
K56 Lg56 Lflux56 1

Cg56 111 0 50.0000fF 
Lg56 111 112 57.0000pH
B56 111 112 10055 jj0 
Cgg56 112 0 50.0000fF
Vmeas56 112 113 0V

*Flux Biasing 
Idc57 0 50057 pwl(0 0uA 5ns 14.0680uA) 
Lflux57 50057 0 57.0000pH 
K57 Lg57 Lflux57 1

Cg57 113 0 50.0000fF 
Lg57 113 114 57.0000pH
B57 113 114 10056 jj0 
Cgg57 114 0 50.0000fF
Vmeas57 114 115 0V

*Flux Biasing 
Idc58 0 50058 pwl(0 0uA 5ns 14.0680uA) 
Lflux58 50058 0 57.0000pH 
K58 Lg58 Lflux58 1

Cg58 115 0 50.0000fF 
Lg58 115 116 57.0000pH
B58 115 116 10057 jj0 
Cgg58 116 0 50.0000fF
Vmeas58 116 117 0V

*Flux Biasing 
Idc59 0 50059 pwl(0 0uA 5ns 14.0680uA) 
Lflux59 50059 0 57.0000pH 
K59 Lg59 Lflux59 1

Cg59 117 0 50.0000fF 
Lg59 117 118 57.0000pH
B59 117 118 10058 jj0 
Cgg59 118 0 50.0000fF
Vmeas59 118 119 0V

*Flux Biasing 
Idc60 0 50060 pwl(0 0uA 5ns 14.0680uA) 
Lflux60 50060 0 57.0000pH 
K60 Lg60 Lflux60 1

Cg60 119 0 50.0000fF 
Lg60 119 120 57.0000pH
B60 119 120 10059 jj0 
Cgg60 120 0 50.0000fF
Vmeas60 120 121 0V

*Flux Biasing 
Idc61 0 50061 pwl(0 0uA 5ns 14.0680uA) 
Lflux61 50061 0 57.0000pH 
K61 Lg61 Lflux61 1

Cg61 121 0 50.0000fF 
Lg61 121 122 57.0000pH
B61 121 122 10060 jj0 
Cgg61 122 0 50.0000fF
Vmeas61 122 123 0V

*Flux Biasing 
Idc62 0 50062 pwl(0 0uA 5ns 14.0680uA) 
Lflux62 50062 0 57.0000pH 
K62 Lg62 Lflux62 1

Cg62 123 0 50.0000fF 
Lg62 123 124 57.0000pH
B62 123 124 10061 jj0 
Cgg62 124 0 50.0000fF
Vmeas62 124 125 0V

*Flux Biasing 
Idc63 0 50063 pwl(0 0uA 5ns 14.0680uA) 
Lflux63 50063 0 57.0000pH 
K63 Lg63 Lflux63 1

Cg63 125 0 50.0000fF 
Lg63 125 126 57.0000pH
B63 125 126 10062 jj0 
Cgg63 126 0 50.0000fF
Vmeas63 126 127 0V

*Flux Biasing 
Idc64 0 50064 pwl(0 0uA 5ns 14.0680uA) 
Lflux64 50064 0 57.0000pH 
K64 Lg64 Lflux64 1

Cg64 127 0 50.0000fF 
Lg64 127 128 57.0000pH
B64 127 128 10063 jj0 
Cgg64 128 0 50.0000fF
Vmeas64 128 129 0V

*Flux Biasing 
Idc65 0 50065 pwl(0 0uA 5ns 14.0680uA) 
Lflux65 50065 0 57.0000pH 
K65 Lg65 Lflux65 1

Cg65 129 0 50.0000fF 
Lg65 129 130 57.0000pH
B65 129 130 10064 jj0 
Cgg65 130 0 50.0000fF
Vmeas65 130 131 0V

*Flux Biasing 
Idc66 0 50066 pwl(0 0uA 5ns 14.0680uA) 
Lflux66 50066 0 57.0000pH 
K66 Lg66 Lflux66 1

Cg66 131 0 50.0000fF 
Lg66 131 132 57.0000pH
B66 131 132 10065 jj0 
Cgg66 132 0 50.0000fF
Vmeas66 132 133 0V

*Flux Biasing 
Idc67 0 50067 pwl(0 0uA 5ns 14.0680uA) 
Lflux67 50067 0 57.0000pH 
K67 Lg67 Lflux67 1

Cg67 133 0 50.0000fF 
Lg67 133 134 57.0000pH
B67 133 134 10066 jj0 
Cgg67 134 0 50.0000fF
Vmeas67 134 135 0V

*Flux Biasing 
Idc68 0 50068 pwl(0 0uA 5ns 14.0680uA) 
Lflux68 50068 0 57.0000pH 
K68 Lg68 Lflux68 1

Cg68 135 0 50.0000fF 
Lg68 135 136 57.0000pH
B68 135 136 10067 jj0 
Cgg68 136 0 50.0000fF
Vmeas68 136 137 0V

*Flux Biasing 
Idc69 0 50069 pwl(0 0uA 5ns 14.0680uA) 
Lflux69 50069 0 57.0000pH 
K69 Lg69 Lflux69 1

Cg69 137 0 50.0000fF 
Lg69 137 138 57.0000pH
B69 137 138 10068 jj0 
Cgg69 138 0 50.0000fF
Vmeas69 138 139 0V

*Flux Biasing 
Idc70 0 50070 pwl(0 0uA 5ns 14.0680uA) 
Lflux70 50070 0 57.0000pH 
K70 Lg70 Lflux70 1

Cg70 139 0 50.0000fF 
Lg70 139 140 57.0000pH
B70 139 140 10069 jj0 
Cgg70 140 0 50.0000fF
Vmeas70 140 141 0V

*Flux Biasing 
Idc71 0 50071 pwl(0 0uA 5ns 14.0680uA) 
Lflux71 50071 0 57.0000pH 
K71 Lg71 Lflux71 1

Cg71 141 0 50.0000fF 
Lg71 141 142 57.0000pH
B71 141 142 10070 jj0 
Cgg71 142 0 50.0000fF
Vmeas71 142 143 0V

*Flux Biasing 
Idc72 0 50072 pwl(0 0uA 5ns 14.0680uA) 
Lflux72 50072 0 57.0000pH 
K72 Lg72 Lflux72 1

Cg72 143 0 50.0000fF 
Lg72 143 144 57.0000pH
B72 143 144 10071 jj0 
Cgg72 144 0 50.0000fF
Vmeas72 144 145 0V

*Flux Biasing 
Idc73 0 50073 pwl(0 0uA 5ns 14.0680uA) 
Lflux73 50073 0 57.0000pH 
K73 Lg73 Lflux73 1

Cg73 145 0 50.0000fF 
Lg73 145 146 57.0000pH
B73 145 146 10072 jj0 
Cgg73 146 0 50.0000fF
Vmeas73 146 147 0V

*Flux Biasing 
Idc74 0 50074 pwl(0 0uA 5ns 14.0680uA) 
Lflux74 50074 0 57.0000pH 
K74 Lg74 Lflux74 1

Cg74 147 0 50.0000fF 
Lg74 147 148 57.0000pH
B74 147 148 10073 jj0 
Cgg74 148 0 50.0000fF
Vmeas74 148 149 0V

*Flux Biasing 
Idc75 0 50075 pwl(0 0uA 5ns 14.0680uA) 
Lflux75 50075 0 57.0000pH 
K75 Lg75 Lflux75 1

Cg75 149 0 50.0000fF 
Lg75 149 150 57.0000pH
B75 149 150 10074 jj0 
Cgg75 150 0 50.0000fF
Vmeas75 150 151 0V

*Flux Biasing 
Idc76 0 50076 pwl(0 0uA 5ns 14.0680uA) 
Lflux76 50076 0 57.0000pH 
K76 Lg76 Lflux76 1

Cg76 151 0 50.0000fF 
Lg76 151 152 57.0000pH
B76 151 152 10075 jj0 
Cgg76 152 0 50.0000fF
Vmeas76 152 153 0V

*Flux Biasing 
Idc77 0 50077 pwl(0 0uA 5ns 14.0680uA) 
Lflux77 50077 0 57.0000pH 
K77 Lg77 Lflux77 1

Cg77 153 0 50.0000fF 
Lg77 153 154 57.0000pH
B77 153 154 10076 jj0 
Cgg77 154 0 50.0000fF
Vmeas77 154 155 0V

*Flux Biasing 
Idc78 0 50078 pwl(0 0uA 5ns 14.0680uA) 
Lflux78 50078 0 57.0000pH 
K78 Lg78 Lflux78 1

Cg78 155 0 50.0000fF 
Lg78 155 156 57.0000pH
B78 155 156 10077 jj0 
Cgg78 156 0 50.0000fF
Vmeas78 156 157 0V

*Flux Biasing 
Idc79 0 50079 pwl(0 0uA 5ns 14.0680uA) 
Lflux79 50079 0 57.0000pH 
K79 Lg79 Lflux79 1

Cg79 157 0 50.0000fF 
Lg79 157 158 57.0000pH
B79 157 158 10078 jj0 
Cgg79 158 0 50.0000fF
Vmeas79 158 159 0V

*Flux Biasing 
Idc80 0 50080 pwl(0 0uA 5ns 14.0680uA) 
Lflux80 50080 0 57.0000pH 
K80 Lg80 Lflux80 1

Cg80 159 0 50.0000fF 
Lg80 159 160 57.0000pH
B80 159 160 10079 jj0 
Cgg80 160 0 50.0000fF
Vmeas80 160 161 0V

*Flux Biasing 
Idc81 0 50081 pwl(0 0uA 5ns 14.0680uA) 
Lflux81 50081 0 57.0000pH 
K81 Lg81 Lflux81 1

Cg81 161 0 50.0000fF 
Lg81 161 162 57.0000pH
B81 161 162 10080 jj0 
Cgg81 162 0 50.0000fF
Vmeas81 162 163 0V

*Flux Biasing 
Idc82 0 50082 pwl(0 0uA 5ns 14.0680uA) 
Lflux82 50082 0 57.0000pH 
K82 Lg82 Lflux82 1

Cg82 163 0 50.0000fF 
Lg82 163 164 57.0000pH
B82 163 164 10081 jj0 
Cgg82 164 0 50.0000fF
Vmeas82 164 165 0V

*Flux Biasing 
Idc83 0 50083 pwl(0 0uA 5ns 14.0680uA) 
Lflux83 50083 0 57.0000pH 
K83 Lg83 Lflux83 1

Cg83 165 0 50.0000fF 
Lg83 165 166 57.0000pH
B83 165 166 10082 jj0 
Cgg83 166 0 50.0000fF
Vmeas83 166 167 0V

*Flux Biasing 
Idc84 0 50084 pwl(0 0uA 5ns 14.0680uA) 
Lflux84 50084 0 57.0000pH 
K84 Lg84 Lflux84 1

Cg84 167 0 50.0000fF 
Lg84 167 168 57.0000pH
B84 167 168 10083 jj0 
Cgg84 168 0 50.0000fF
Vmeas84 168 169 0V

*Flux Biasing 
Idc85 0 50085 pwl(0 0uA 5ns 14.0680uA) 
Lflux85 50085 0 57.0000pH 
K85 Lg85 Lflux85 1

Cg85 169 0 50.0000fF 
Lg85 169 170 57.0000pH
B85 169 170 10084 jj0 
Cgg85 170 0 50.0000fF
Vmeas85 170 171 0V

*Flux Biasing 
Idc86 0 50086 pwl(0 0uA 5ns 14.0680uA) 
Lflux86 50086 0 57.0000pH 
K86 Lg86 Lflux86 1

Cg86 171 0 50.0000fF 
Lg86 171 172 57.0000pH
B86 171 172 10085 jj0 
Cgg86 172 0 50.0000fF
Vmeas86 172 173 0V

*Flux Biasing 
Idc87 0 50087 pwl(0 0uA 5ns 14.0680uA) 
Lflux87 50087 0 57.0000pH 
K87 Lg87 Lflux87 1

Cg87 173 0 50.0000fF 
Lg87 173 174 57.0000pH
B87 173 174 10086 jj0 
Cgg87 174 0 50.0000fF
Vmeas87 174 175 0V

*Flux Biasing 
Idc88 0 50088 pwl(0 0uA 5ns 14.0680uA) 
Lflux88 50088 0 57.0000pH 
K88 Lg88 Lflux88 1

Cg88 175 0 50.0000fF 
Lg88 175 176 57.0000pH
B88 175 176 10087 jj0 
Cgg88 176 0 50.0000fF
Vmeas88 176 177 0V

*Flux Biasing 
Idc89 0 50089 pwl(0 0uA 5ns 14.0680uA) 
Lflux89 50089 0 57.0000pH 
K89 Lg89 Lflux89 1

Cg89 177 0 50.0000fF 
Lg89 177 178 57.0000pH
B89 177 178 10088 jj0 
Cgg89 178 0 50.0000fF
Vmeas89 178 179 0V

*Flux Biasing 
Idc90 0 50090 pwl(0 0uA 5ns 14.0680uA) 
Lflux90 50090 0 57.0000pH 
K90 Lg90 Lflux90 1

Cg90 179 0 50.0000fF 
Lg90 179 180 57.0000pH
B90 179 180 10089 jj0 
Cgg90 180 0 50.0000fF
Vmeas90 180 181 0V

*Flux Biasing 
Idc91 0 50091 pwl(0 0uA 5ns 14.0680uA) 
Lflux91 50091 0 57.0000pH 
K91 Lg91 Lflux91 1

Cg91 181 0 50.0000fF 
Lg91 181 182 57.0000pH
B91 181 182 10090 jj0 
Cgg91 182 0 50.0000fF
Vmeas91 182 183 0V

*Flux Biasing 
Idc92 0 50092 pwl(0 0uA 5ns 14.0680uA) 
Lflux92 50092 0 57.0000pH 
K92 Lg92 Lflux92 1

Cg92 183 0 50.0000fF 
Lg92 183 184 57.0000pH
B92 183 184 10091 jj0 
Cgg92 184 0 50.0000fF
Vmeas92 184 185 0V

*Flux Biasing 
Idc93 0 50093 pwl(0 0uA 5ns 14.0680uA) 
Lflux93 50093 0 57.0000pH 
K93 Lg93 Lflux93 1

Cg93 185 0 50.0000fF 
Lg93 185 186 57.0000pH
B93 185 186 10092 jj0 
Cgg93 186 0 50.0000fF
Vmeas93 186 187 0V

*Flux Biasing 
Idc94 0 50094 pwl(0 0uA 5ns 14.0680uA) 
Lflux94 50094 0 57.0000pH 
K94 Lg94 Lflux94 1

Cg94 187 0 50.0000fF 
Lg94 187 188 57.0000pH
B94 187 188 10093 jj0 
Cgg94 188 0 50.0000fF
Vmeas94 188 189 0V

*Flux Biasing 
Idc95 0 50095 pwl(0 0uA 5ns 14.0680uA) 
Lflux95 50095 0 57.0000pH 
K95 Lg95 Lflux95 1

Cg95 189 0 50.0000fF 
Lg95 189 190 57.0000pH
B95 189 190 10094 jj0 
Cgg95 190 0 50.0000fF
Vmeas95 190 191 0V

*Flux Biasing 
Idc96 0 50096 pwl(0 0uA 5ns 14.0680uA) 
Lflux96 50096 0 57.0000pH 
K96 Lg96 Lflux96 1

Cg96 191 0 50.0000fF 
Lg96 191 192 57.0000pH
B96 191 192 10095 jj0 
Cgg96 192 0 50.0000fF
Vmeas96 192 193 0V

*Flux Biasing 
Idc97 0 50097 pwl(0 0uA 5ns 14.0680uA) 
Lflux97 50097 0 57.0000pH 
K97 Lg97 Lflux97 1

Cg97 193 0 50.0000fF 
Lg97 193 194 57.0000pH
B97 193 194 10096 jj0 
Cgg97 194 0 50.0000fF
Vmeas97 194 195 0V

*Flux Biasing 
Idc98 0 50098 pwl(0 0uA 5ns 14.0680uA) 
Lflux98 50098 0 57.0000pH 
K98 Lg98 Lflux98 1

Cg98 195 0 50.0000fF 
Lg98 195 196 57.0000pH
B98 195 196 10097 jj0 
Cgg98 196 0 50.0000fF
Vmeas98 196 197 0V

*Flux Biasing 
Idc99 0 50099 pwl(0 0uA 5ns 14.0680uA) 
Lflux99 50099 0 57.0000pH 
K99 Lg99 Lflux99 1

Cg99 197 0 50.0000fF 
Lg99 197 198 57.0000pH
B99 197 198 10098 jj0 
Cgg99 198 0 50.0000fF
Vmeas99 198 199 0V

*Flux Biasing 
Idc100 0 50100 pwl(0 0uA 5ns 14.0680uA) 
Lflux100 50100 0 57.0000pH 
K100 Lg100 Lflux100 1

Cg100 199 0 50.0000fF 
Lg100 199 200 57.0000pH
B100 199 200 10099 jj0 
Cgg100 200 0 50.0000fF
Vmeas100 200 201 0V

*Flux Biasing 
Idc101 0 50101 pwl(0 0uA 5ns 14.0680uA) 
Lflux101 50101 0 57.0000pH 
K101 Lg101 Lflux101 1

Cg101 201 0 50.0000fF 
Lg101 201 202 57.0000pH
B101 201 202 10100 jj0 
Cgg101 202 0 50.0000fF
Vmeas101 202 203 0V

*Flux Biasing 
Idc102 0 50102 pwl(0 0uA 5ns 14.0680uA) 
Lflux102 50102 0 57.0000pH 
K102 Lg102 Lflux102 1

Cg102 203 0 50.0000fF 
Lg102 203 204 57.0000pH
B102 203 204 10101 jj0 
Cgg102 204 0 50.0000fF
Vmeas102 204 205 0V

*Flux Biasing 
Idc103 0 50103 pwl(0 0uA 5ns 14.0680uA) 
Lflux103 50103 0 57.0000pH 
K103 Lg103 Lflux103 1

Cg103 205 0 50.0000fF 
Lg103 205 206 57.0000pH
B103 205 206 10102 jj0 
Cgg103 206 0 50.0000fF
Vmeas103 206 207 0V

*Flux Biasing 
Idc104 0 50104 pwl(0 0uA 5ns 14.0680uA) 
Lflux104 50104 0 57.0000pH 
K104 Lg104 Lflux104 1

Cg104 207 0 50.0000fF 
Lg104 207 208 57.0000pH
B104 207 208 10103 jj0 
Cgg104 208 0 50.0000fF
Vmeas104 208 209 0V

*Flux Biasing 
Idc105 0 50105 pwl(0 0uA 5ns 14.0680uA) 
Lflux105 50105 0 57.0000pH 
K105 Lg105 Lflux105 1

Cg105 209 0 50.0000fF 
Lg105 209 210 57.0000pH
B105 209 210 10104 jj0 
Cgg105 210 0 50.0000fF
Vmeas105 210 211 0V

*Flux Biasing 
Idc106 0 50106 pwl(0 0uA 5ns 14.0680uA) 
Lflux106 50106 0 57.0000pH 
K106 Lg106 Lflux106 1

Cg106 211 0 50.0000fF 
Lg106 211 212 57.0000pH
B106 211 212 10105 jj0 
Cgg106 212 0 50.0000fF
Vmeas106 212 213 0V

*Flux Biasing 
Idc107 0 50107 pwl(0 0uA 5ns 14.0680uA) 
Lflux107 50107 0 57.0000pH 
K107 Lg107 Lflux107 1

Cg107 213 0 50.0000fF 
Lg107 213 214 57.0000pH
B107 213 214 10106 jj0 
Cgg107 214 0 50.0000fF
Vmeas107 214 215 0V

*Flux Biasing 
Idc108 0 50108 pwl(0 0uA 5ns 14.0680uA) 
Lflux108 50108 0 57.0000pH 
K108 Lg108 Lflux108 1

Cg108 215 0 50.0000fF 
Lg108 215 216 57.0000pH
B108 215 216 10107 jj0 
Cgg108 216 0 50.0000fF
Vmeas108 216 217 0V

*Flux Biasing 
Idc109 0 50109 pwl(0 0uA 5ns 14.0680uA) 
Lflux109 50109 0 57.0000pH 
K109 Lg109 Lflux109 1

Cg109 217 0 50.0000fF 
Lg109 217 218 57.0000pH
B109 217 218 10108 jj0 
Cgg109 218 0 50.0000fF
Vmeas109 218 219 0V

*Flux Biasing 
Idc110 0 50110 pwl(0 0uA 5ns 14.0680uA) 
Lflux110 50110 0 57.0000pH 
K110 Lg110 Lflux110 1

Cg110 219 0 50.0000fF 
Lg110 219 220 57.0000pH
B110 219 220 10109 jj0 
Cgg110 220 0 50.0000fF
Vmeas110 220 221 0V

*Flux Biasing 
Idc111 0 50111 pwl(0 0uA 5ns 14.0680uA) 
Lflux111 50111 0 57.0000pH 
K111 Lg111 Lflux111 1

Cg111 221 0 50.0000fF 
Lg111 221 222 57.0000pH
B111 221 222 10110 jj0 
Cgg111 222 0 50.0000fF
Vmeas111 222 223 0V

*Flux Biasing 
Idc112 0 50112 pwl(0 0uA 5ns 14.0680uA) 
Lflux112 50112 0 57.0000pH 
K112 Lg112 Lflux112 1

Cg112 223 0 50.0000fF 
Lg112 223 224 57.0000pH
B112 223 224 10111 jj0 
Cgg112 224 0 50.0000fF
Vmeas112 224 225 0V

*Flux Biasing 
Idc113 0 50113 pwl(0 0uA 5ns 14.0680uA) 
Lflux113 50113 0 57.0000pH 
K113 Lg113 Lflux113 1

Cg113 225 0 50.0000fF 
Lg113 225 226 57.0000pH
B113 225 226 10112 jj0 
Cgg113 226 0 50.0000fF
Vmeas113 226 227 0V

*Flux Biasing 
Idc114 0 50114 pwl(0 0uA 5ns 14.0680uA) 
Lflux114 50114 0 57.0000pH 
K114 Lg114 Lflux114 1

Cg114 227 0 50.0000fF 
Lg114 227 228 57.0000pH
B114 227 228 10113 jj0 
Cgg114 228 0 50.0000fF
Vmeas114 228 229 0V

*Flux Biasing 
Idc115 0 50115 pwl(0 0uA 5ns 14.0680uA) 
Lflux115 50115 0 57.0000pH 
K115 Lg115 Lflux115 1

Cg115 229 0 50.0000fF 
Lg115 229 230 57.0000pH
B115 229 230 10114 jj0 
Cgg115 230 0 50.0000fF
Vmeas115 230 231 0V

*Flux Biasing 
Idc116 0 50116 pwl(0 0uA 5ns 14.0680uA) 
Lflux116 50116 0 57.0000pH 
K116 Lg116 Lflux116 1

Cg116 231 0 50.0000fF 
Lg116 231 232 57.0000pH
B116 231 232 10115 jj0 
Cgg116 232 0 50.0000fF
Vmeas116 232 233 0V

*Flux Biasing 
Idc117 0 50117 pwl(0 0uA 5ns 14.0680uA) 
Lflux117 50117 0 57.0000pH 
K117 Lg117 Lflux117 1

Cg117 233 0 50.0000fF 
Lg117 233 234 57.0000pH
B117 233 234 10116 jj0 
Cgg117 234 0 50.0000fF
Vmeas117 234 235 0V

*Flux Biasing 
Idc118 0 50118 pwl(0 0uA 5ns 14.0680uA) 
Lflux118 50118 0 57.0000pH 
K118 Lg118 Lflux118 1

Cg118 235 0 50.0000fF 
Lg118 235 236 57.0000pH
B118 235 236 10117 jj0 
Cgg118 236 0 50.0000fF
Vmeas118 236 237 0V

*Flux Biasing 
Idc119 0 50119 pwl(0 0uA 5ns 14.0680uA) 
Lflux119 50119 0 57.0000pH 
K119 Lg119 Lflux119 1

Cg119 237 0 50.0000fF 
Lg119 237 238 57.0000pH
B119 237 238 10118 jj0 
Cgg119 238 0 50.0000fF
Vmeas119 238 239 0V

*Flux Biasing 
Idc120 0 50120 pwl(0 0uA 5ns 14.0680uA) 
Lflux120 50120 0 57.0000pH 
K120 Lg120 Lflux120 1

Cg120 239 0 50.0000fF 
Lg120 239 240 57.0000pH
B120 239 240 10119 jj0 
Cgg120 240 0 50.0000fF
Vmeas120 240 241 0V

*Flux Biasing 
Idc121 0 50121 pwl(0 0uA 5ns 14.0680uA) 
Lflux121 50121 0 57.0000pH 
K121 Lg121 Lflux121 1

Cg121 241 0 50.0000fF 
Lg121 241 242 57.0000pH
B121 241 242 10120 jj0 
Cgg121 242 0 50.0000fF
Vmeas121 242 243 0V

*Flux Biasing 
Idc122 0 50122 pwl(0 0uA 5ns 14.0680uA) 
Lflux122 50122 0 57.0000pH 
K122 Lg122 Lflux122 1

Cg122 243 0 50.0000fF 
Lg122 243 244 57.0000pH
B122 243 244 10121 jj0 
Cgg122 244 0 50.0000fF
Vmeas122 244 245 0V

*Flux Biasing 
Idc123 0 50123 pwl(0 0uA 5ns 14.0680uA) 
Lflux123 50123 0 57.0000pH 
K123 Lg123 Lflux123 1

Cg123 245 0 50.0000fF 
Lg123 245 246 57.0000pH
B123 245 246 10122 jj0 
Cgg123 246 0 50.0000fF
Vmeas123 246 247 0V

*Flux Biasing 
Idc124 0 50124 pwl(0 0uA 5ns 14.0680uA) 
Lflux124 50124 0 57.0000pH 
K124 Lg124 Lflux124 1

Cg124 247 0 50.0000fF 
Lg124 247 248 57.0000pH
B124 247 248 10123 jj0 
Cgg124 248 0 50.0000fF
Vmeas124 248 249 0V

*Flux Biasing 
Idc125 0 50125 pwl(0 0uA 5ns 14.0680uA) 
Lflux125 50125 0 57.0000pH 
K125 Lg125 Lflux125 1

Cg125 249 0 50.0000fF 
Lg125 249 250 57.0000pH
B125 249 250 10124 jj0 
Cgg125 250 0 50.0000fF
Vmeas125 250 251 0V

*Flux Biasing 
Idc126 0 50126 pwl(0 0uA 5ns 14.0680uA) 
Lflux126 50126 0 57.0000pH 
K126 Lg126 Lflux126 1

Cg126 251 0 50.0000fF 
Lg126 251 252 57.0000pH
B126 251 252 10125 jj0 
Cgg126 252 0 50.0000fF
Vmeas126 252 253 0V

*Flux Biasing 
Idc127 0 50127 pwl(0 0uA 5ns 14.0680uA) 
Lflux127 50127 0 57.0000pH 
K127 Lg127 Lflux127 1

Cg127 253 0 50.0000fF 
Lg127 253 254 57.0000pH
B127 253 254 10126 jj0 
Cgg127 254 0 50.0000fF
Vmeas127 254 255 0V

*Flux Biasing 
Idc128 0 50128 pwl(0 0uA 5ns 14.0680uA) 
Lflux128 50128 0 57.0000pH 
K128 Lg128 Lflux128 1

Cg128 255 0 50.0000fF 
Lg128 255 256 57.0000pH
B128 255 256 10127 jj0 
Cgg128 256 0 50.0000fF
Vmeas128 256 257 0V

*Flux Biasing 
Idc129 0 50129 pwl(0 0uA 5ns 14.0680uA) 
Lflux129 50129 0 57.0000pH 
K129 Lg129 Lflux129 1

Cg129 257 0 50.0000fF 
Lg129 257 258 57.0000pH
B129 257 258 10128 jj0 
Cgg129 258 0 50.0000fF
Vmeas129 258 259 0V

*Flux Biasing 
Idc130 0 50130 pwl(0 0uA 5ns 14.0680uA) 
Lflux130 50130 0 57.0000pH 
K130 Lg130 Lflux130 1

Cg130 259 0 50.0000fF 
Lg130 259 260 57.0000pH
B130 259 260 10129 jj0 
Cgg130 260 0 50.0000fF
Vmeas130 260 261 0V

*Flux Biasing 
Idc131 0 50131 pwl(0 0uA 5ns 14.0680uA) 
Lflux131 50131 0 57.0000pH 
K131 Lg131 Lflux131 1

Cg131 261 0 50.0000fF 
Lg131 261 262 57.0000pH
B131 261 262 10130 jj0 
Cgg131 262 0 50.0000fF
Vmeas131 262 263 0V

*Flux Biasing 
Idc132 0 50132 pwl(0 0uA 5ns 14.0680uA) 
Lflux132 50132 0 57.0000pH 
K132 Lg132 Lflux132 1

Cg132 263 0 50.0000fF 
Lg132 263 264 57.0000pH
B132 263 264 10131 jj0 
Cgg132 264 0 50.0000fF
Vmeas132 264 265 0V

*Flux Biasing 
Idc133 0 50133 pwl(0 0uA 5ns 14.0680uA) 
Lflux133 50133 0 57.0000pH 
K133 Lg133 Lflux133 1

Cg133 265 0 50.0000fF 
Lg133 265 266 57.0000pH
B133 265 266 10132 jj0 
Cgg133 266 0 50.0000fF
Vmeas133 266 267 0V

*Flux Biasing 
Idc134 0 50134 pwl(0 0uA 5ns 14.0680uA) 
Lflux134 50134 0 57.0000pH 
K134 Lg134 Lflux134 1

Cg134 267 0 50.0000fF 
Lg134 267 268 57.0000pH
B134 267 268 10133 jj0 
Cgg134 268 0 50.0000fF
Vmeas134 268 269 0V

*Flux Biasing 
Idc135 0 50135 pwl(0 0uA 5ns 14.0680uA) 
Lflux135 50135 0 57.0000pH 
K135 Lg135 Lflux135 1

Cg135 269 0 50.0000fF 
Lg135 269 270 57.0000pH
B135 269 270 10134 jj0 
Cgg135 270 0 50.0000fF
Vmeas135 270 271 0V

*Flux Biasing 
Idc136 0 50136 pwl(0 0uA 5ns 14.0680uA) 
Lflux136 50136 0 57.0000pH 
K136 Lg136 Lflux136 1

Cg136 271 0 50.0000fF 
Lg136 271 272 57.0000pH
B136 271 272 10135 jj0 
Cgg136 272 0 50.0000fF
Vmeas136 272 273 0V

*Flux Biasing 
Idc137 0 50137 pwl(0 0uA 5ns 14.0680uA) 
Lflux137 50137 0 57.0000pH 
K137 Lg137 Lflux137 1

Cg137 273 0 50.0000fF 
Lg137 273 274 57.0000pH
B137 273 274 10136 jj0 
Cgg137 274 0 50.0000fF
Vmeas137 274 275 0V

*Flux Biasing 
Idc138 0 50138 pwl(0 0uA 5ns 14.0680uA) 
Lflux138 50138 0 57.0000pH 
K138 Lg138 Lflux138 1

Cg138 275 0 50.0000fF 
Lg138 275 276 57.0000pH
B138 275 276 10137 jj0 
Cgg138 276 0 50.0000fF
Vmeas138 276 277 0V

*Flux Biasing 
Idc139 0 50139 pwl(0 0uA 5ns 14.0680uA) 
Lflux139 50139 0 57.0000pH 
K139 Lg139 Lflux139 1

Cg139 277 0 50.0000fF 
Lg139 277 278 57.0000pH
B139 277 278 10138 jj0 
Cgg139 278 0 50.0000fF
Vmeas139 278 279 0V

*Flux Biasing 
Idc140 0 50140 pwl(0 0uA 5ns 14.0680uA) 
Lflux140 50140 0 57.0000pH 
K140 Lg140 Lflux140 1

Cg140 279 0 50.0000fF 
Lg140 279 280 57.0000pH
B140 279 280 10139 jj0 
Cgg140 280 0 50.0000fF
Vmeas140 280 281 0V

*Flux Biasing 
Idc141 0 50141 pwl(0 0uA 5ns 14.0680uA) 
Lflux141 50141 0 57.0000pH 
K141 Lg141 Lflux141 1

Cg141 281 0 50.0000fF 
Lg141 281 282 57.0000pH
B141 281 282 10140 jj0 
Cgg141 282 0 50.0000fF
Vmeas141 282 283 0V

*Flux Biasing 
Idc142 0 50142 pwl(0 0uA 5ns 14.0680uA) 
Lflux142 50142 0 57.0000pH 
K142 Lg142 Lflux142 1

Cg142 283 0 50.0000fF 
Lg142 283 284 57.0000pH
B142 283 284 10141 jj0 
Cgg142 284 0 50.0000fF
Vmeas142 284 285 0V

*Flux Biasing 
Idc143 0 50143 pwl(0 0uA 5ns 14.0680uA) 
Lflux143 50143 0 57.0000pH 
K143 Lg143 Lflux143 1

Cg143 285 0 50.0000fF 
Lg143 285 286 57.0000pH
B143 285 286 10142 jj0 
Cgg143 286 0 50.0000fF
Vmeas143 286 287 0V

*Flux Biasing 
Idc144 0 50144 pwl(0 0uA 5ns 14.0680uA) 
Lflux144 50144 0 57.0000pH 
K144 Lg144 Lflux144 1

Cg144 287 0 50.0000fF 
Lg144 287 288 57.0000pH
B144 287 288 10143 jj0 
Cgg144 288 0 50.0000fF
Vmeas144 288 289 0V

*Flux Biasing 
Idc145 0 50145 pwl(0 0uA 5ns 14.0680uA) 
Lflux145 50145 0 57.0000pH 
K145 Lg145 Lflux145 1

Cg145 289 0 50.0000fF 
Lg145 289 290 57.0000pH
B145 289 290 10144 jj0 
Cgg145 290 0 50.0000fF
Vmeas145 290 291 0V

*Flux Biasing 
Idc146 0 50146 pwl(0 0uA 5ns 14.0680uA) 
Lflux146 50146 0 57.0000pH 
K146 Lg146 Lflux146 1

Cg146 291 0 50.0000fF 
Lg146 291 292 57.0000pH
B146 291 292 10145 jj0 
Cgg146 292 0 50.0000fF
Vmeas146 292 293 0V

*Flux Biasing 
Idc147 0 50147 pwl(0 0uA 5ns 14.0680uA) 
Lflux147 50147 0 57.0000pH 
K147 Lg147 Lflux147 1

Cg147 293 0 50.0000fF 
Lg147 293 294 57.0000pH
B147 293 294 10146 jj0 
Cgg147 294 0 50.0000fF
Vmeas147 294 295 0V

*Flux Biasing 
Idc148 0 50148 pwl(0 0uA 5ns 14.0680uA) 
Lflux148 50148 0 57.0000pH 
K148 Lg148 Lflux148 1

Cg148 295 0 50.0000fF 
Lg148 295 296 57.0000pH
B148 295 296 10147 jj0 
Cgg148 296 0 50.0000fF
Vmeas148 296 297 0V

*Flux Biasing 
Idc149 0 50149 pwl(0 0uA 5ns 14.0680uA) 
Lflux149 50149 0 57.0000pH 
K149 Lg149 Lflux149 1

Cg149 297 0 50.0000fF 
Lg149 297 298 57.0000pH
B149 297 298 10148 jj0 
Cgg149 298 0 50.0000fF
Vmeas149 298 299 0V

*Flux Biasing 
Idc150 0 50150 pwl(0 0uA 5ns 14.0680uA) 
Lflux150 50150 0 57.0000pH 
K150 Lg150 Lflux150 1

Cg150 299 0 50.0000fF 
Lg150 299 300 57.0000pH
B150 299 300 10149 jj0 
Cgg150 300 0 50.0000fF
Vmeas150 300 301 0V

*Flux Biasing 
Idc151 0 50151 pwl(0 0uA 5ns 14.0680uA) 
Lflux151 50151 0 57.0000pH 
K151 Lg151 Lflux151 1

Cg151 301 0 50.0000fF 
Lg151 301 302 57.0000pH
B151 301 302 10150 jj0 
Cgg151 302 0 50.0000fF
Vmeas151 302 303 0V

*Flux Biasing 
Idc152 0 50152 pwl(0 0uA 5ns 14.0680uA) 
Lflux152 50152 0 57.0000pH 
K152 Lg152 Lflux152 1

Cg152 303 0 50.0000fF 
Lg152 303 304 57.0000pH
B152 303 304 10151 jj0 
Cgg152 304 0 50.0000fF
Vmeas152 304 305 0V

*Flux Biasing 
Idc153 0 50153 pwl(0 0uA 5ns 14.0680uA) 
Lflux153 50153 0 57.0000pH 
K153 Lg153 Lflux153 1

Cg153 305 0 50.0000fF 
Lg153 305 306 57.0000pH
B153 305 306 10152 jj0 
Cgg153 306 0 50.0000fF
Vmeas153 306 307 0V

*Flux Biasing 
Idc154 0 50154 pwl(0 0uA 5ns 14.0680uA) 
Lflux154 50154 0 57.0000pH 
K154 Lg154 Lflux154 1

Cg154 307 0 50.0000fF 
Lg154 307 308 57.0000pH
B154 307 308 10153 jj0 
Cgg154 308 0 50.0000fF
Vmeas154 308 309 0V

*Flux Biasing 
Idc155 0 50155 pwl(0 0uA 5ns 14.0680uA) 
Lflux155 50155 0 57.0000pH 
K155 Lg155 Lflux155 1

Cg155 309 0 50.0000fF 
Lg155 309 310 57.0000pH
B155 309 310 10154 jj0 
Cgg155 310 0 50.0000fF
Vmeas155 310 311 0V

*Flux Biasing 
Idc156 0 50156 pwl(0 0uA 5ns 14.0680uA) 
Lflux156 50156 0 57.0000pH 
K156 Lg156 Lflux156 1

Cg156 311 0 50.0000fF 
Lg156 311 312 57.0000pH
B156 311 312 10155 jj0 
Cgg156 312 0 50.0000fF
Vmeas156 312 313 0V

*Flux Biasing 
Idc157 0 50157 pwl(0 0uA 5ns 14.0680uA) 
Lflux157 50157 0 57.0000pH 
K157 Lg157 Lflux157 1

Cg157 313 0 50.0000fF 
Lg157 313 314 57.0000pH
B157 313 314 10156 jj0 
Cgg157 314 0 50.0000fF
Vmeas157 314 315 0V

*Flux Biasing 
Idc158 0 50158 pwl(0 0uA 5ns 14.0680uA) 
Lflux158 50158 0 57.0000pH 
K158 Lg158 Lflux158 1

Cg158 315 0 50.0000fF 
Lg158 315 316 57.0000pH
B158 315 316 10157 jj0 
Cgg158 316 0 50.0000fF
Vmeas158 316 317 0V

*Flux Biasing 
Idc159 0 50159 pwl(0 0uA 5ns 14.0680uA) 
Lflux159 50159 0 57.0000pH 
K159 Lg159 Lflux159 1

Cg159 317 0 50.0000fF 
Lg159 317 318 57.0000pH
B159 317 318 10158 jj0 
Cgg159 318 0 50.0000fF
Vmeas159 318 319 0V

*Flux Biasing 
Idc160 0 50160 pwl(0 0uA 5ns 14.0680uA) 
Lflux160 50160 0 57.0000pH 
K160 Lg160 Lflux160 1

Cg160 319 0 50.0000fF 
Lg160 319 320 57.0000pH
B160 319 320 10159 jj0 
Cgg160 320 0 50.0000fF
Vmeas160 320 321 0V

*Flux Biasing 
Idc161 0 50161 pwl(0 0uA 5ns 14.0680uA) 
Lflux161 50161 0 57.0000pH 
K161 Lg161 Lflux161 1

Cg161 321 0 50.0000fF 
Lg161 321 322 57.0000pH
B161 321 322 10160 jj0 
Cgg161 322 0 50.0000fF
Vmeas161 322 323 0V

*Flux Biasing 
Idc162 0 50162 pwl(0 0uA 5ns 14.0680uA) 
Lflux162 50162 0 57.0000pH 
K162 Lg162 Lflux162 1

Cg162 323 0 50.0000fF 
Lg162 323 324 57.0000pH
B162 323 324 10161 jj0 
Cgg162 324 0 50.0000fF
Vmeas162 324 325 0V

*Flux Biasing 
Idc163 0 50163 pwl(0 0uA 5ns 14.0680uA) 
Lflux163 50163 0 57.0000pH 
K163 Lg163 Lflux163 1

Cg163 325 0 50.0000fF 
Lg163 325 326 57.0000pH
B163 325 326 10162 jj0 
Cgg163 326 0 50.0000fF
Vmeas163 326 327 0V

*Flux Biasing 
Idc164 0 50164 pwl(0 0uA 5ns 14.0680uA) 
Lflux164 50164 0 57.0000pH 
K164 Lg164 Lflux164 1

Cg164 327 0 50.0000fF 
Lg164 327 328 57.0000pH
B164 327 328 10163 jj0 
Cgg164 328 0 50.0000fF
Vmeas164 328 329 0V

*Flux Biasing 
Idc165 0 50165 pwl(0 0uA 5ns 14.0680uA) 
Lflux165 50165 0 57.0000pH 
K165 Lg165 Lflux165 1

Cg165 329 0 50.0000fF 
Lg165 329 330 57.0000pH
B165 329 330 10164 jj0 
Cgg165 330 0 50.0000fF
Vmeas165 330 331 0V

*Flux Biasing 
Idc166 0 50166 pwl(0 0uA 5ns 14.0680uA) 
Lflux166 50166 0 57.0000pH 
K166 Lg166 Lflux166 1

Cg166 331 0 50.0000fF 
Lg166 331 332 57.0000pH
B166 331 332 10165 jj0 
Cgg166 332 0 50.0000fF
Vmeas166 332 333 0V

*Flux Biasing 
Idc167 0 50167 pwl(0 0uA 5ns 14.0680uA) 
Lflux167 50167 0 57.0000pH 
K167 Lg167 Lflux167 1

Cg167 333 0 50.0000fF 
Lg167 333 334 57.0000pH
B167 333 334 10166 jj0 
Cgg167 334 0 50.0000fF
Vmeas167 334 335 0V

*Flux Biasing 
Idc168 0 50168 pwl(0 0uA 5ns 14.0680uA) 
Lflux168 50168 0 57.0000pH 
K168 Lg168 Lflux168 1

Cg168 335 0 50.0000fF 
Lg168 335 336 57.0000pH
B168 335 336 10167 jj0 
Cgg168 336 0 50.0000fF
Vmeas168 336 337 0V

*Flux Biasing 
Idc169 0 50169 pwl(0 0uA 5ns 14.0680uA) 
Lflux169 50169 0 57.0000pH 
K169 Lg169 Lflux169 1

Cg169 337 0 50.0000fF 
Lg169 337 338 57.0000pH
B169 337 338 10168 jj0 
Cgg169 338 0 50.0000fF
Vmeas169 338 339 0V

*Flux Biasing 
Idc170 0 50170 pwl(0 0uA 5ns 14.0680uA) 
Lflux170 50170 0 57.0000pH 
K170 Lg170 Lflux170 1

Cg170 339 0 50.0000fF 
Lg170 339 340 57.0000pH
B170 339 340 10169 jj0 
Cgg170 340 0 50.0000fF
Vmeas170 340 341 0V

*Flux Biasing 
Idc171 0 50171 pwl(0 0uA 5ns 14.0680uA) 
Lflux171 50171 0 57.0000pH 
K171 Lg171 Lflux171 1

Cg171 341 0 50.0000fF 
Lg171 341 342 57.0000pH
B171 341 342 10170 jj0 
Cgg171 342 0 50.0000fF
Vmeas171 342 343 0V

*Flux Biasing 
Idc172 0 50172 pwl(0 0uA 5ns 14.0680uA) 
Lflux172 50172 0 57.0000pH 
K172 Lg172 Lflux172 1

Cg172 343 0 50.0000fF 
Lg172 343 344 57.0000pH
B172 343 344 10171 jj0 
Cgg172 344 0 50.0000fF
Vmeas172 344 345 0V

*Flux Biasing 
Idc173 0 50173 pwl(0 0uA 5ns 14.0680uA) 
Lflux173 50173 0 57.0000pH 
K173 Lg173 Lflux173 1

Cg173 345 0 50.0000fF 
Lg173 345 346 57.0000pH
B173 345 346 10172 jj0 
Cgg173 346 0 50.0000fF
Vmeas173 346 347 0V

*Flux Biasing 
Idc174 0 50174 pwl(0 0uA 5ns 14.0680uA) 
Lflux174 50174 0 57.0000pH 
K174 Lg174 Lflux174 1

Cg174 347 0 50.0000fF 
Lg174 347 348 57.0000pH
B174 347 348 10173 jj0 
Cgg174 348 0 50.0000fF
Vmeas174 348 349 0V

*Flux Biasing 
Idc175 0 50175 pwl(0 0uA 5ns 14.0680uA) 
Lflux175 50175 0 57.0000pH 
K175 Lg175 Lflux175 1

Cg175 349 0 50.0000fF 
Lg175 349 350 57.0000pH
B175 349 350 10174 jj0 
Cgg175 350 0 50.0000fF
Vmeas175 350 351 0V

*Flux Biasing 
Idc176 0 50176 pwl(0 0uA 5ns 14.0680uA) 
Lflux176 50176 0 57.0000pH 
K176 Lg176 Lflux176 1

Cg176 351 0 50.0000fF 
Lg176 351 352 57.0000pH
B176 351 352 10175 jj0 
Cgg176 352 0 50.0000fF
Vmeas176 352 353 0V

*Flux Biasing 
Idc177 0 50177 pwl(0 0uA 5ns 14.0680uA) 
Lflux177 50177 0 57.0000pH 
K177 Lg177 Lflux177 1

Cg177 353 0 50.0000fF 
Lg177 353 354 57.0000pH
B177 353 354 10176 jj0 
Cgg177 354 0 50.0000fF
Vmeas177 354 355 0V

*Flux Biasing 
Idc178 0 50178 pwl(0 0uA 5ns 14.0680uA) 
Lflux178 50178 0 57.0000pH 
K178 Lg178 Lflux178 1

Cg178 355 0 50.0000fF 
Lg178 355 356 57.0000pH
B178 355 356 10177 jj0 
Cgg178 356 0 50.0000fF
Vmeas178 356 357 0V

*Flux Biasing 
Idc179 0 50179 pwl(0 0uA 5ns 14.0680uA) 
Lflux179 50179 0 57.0000pH 
K179 Lg179 Lflux179 1

Cg179 357 0 50.0000fF 
Lg179 357 358 57.0000pH
B179 357 358 10178 jj0 
Cgg179 358 0 50.0000fF
Vmeas179 358 359 0V

*Flux Biasing 
Idc180 0 50180 pwl(0 0uA 5ns 14.0680uA) 
Lflux180 50180 0 57.0000pH 
K180 Lg180 Lflux180 1

Cg180 359 0 50.0000fF 
Lg180 359 360 57.0000pH
B180 359 360 10179 jj0 
Cgg180 360 0 50.0000fF
Vmeas180 360 361 0V

*Flux Biasing 
Idc181 0 50181 pwl(0 0uA 5ns 14.0680uA) 
Lflux181 50181 0 57.0000pH 
K181 Lg181 Lflux181 1

Cg181 361 0 50.0000fF 
Lg181 361 362 57.0000pH
B181 361 362 10180 jj0 
Cgg181 362 0 50.0000fF
Vmeas181 362 363 0V

*Flux Biasing 
Idc182 0 50182 pwl(0 0uA 5ns 14.0680uA) 
Lflux182 50182 0 57.0000pH 
K182 Lg182 Lflux182 1

Cg182 363 0 50.0000fF 
Lg182 363 364 57.0000pH
B182 363 364 10181 jj0 
Cgg182 364 0 50.0000fF
Vmeas182 364 365 0V

*Flux Biasing 
Idc183 0 50183 pwl(0 0uA 5ns 14.0680uA) 
Lflux183 50183 0 57.0000pH 
K183 Lg183 Lflux183 1

Cg183 365 0 50.0000fF 
Lg183 365 366 57.0000pH
B183 365 366 10182 jj0 
Cgg183 366 0 50.0000fF
Vmeas183 366 367 0V

*Flux Biasing 
Idc184 0 50184 pwl(0 0uA 5ns 14.0680uA) 
Lflux184 50184 0 57.0000pH 
K184 Lg184 Lflux184 1

Cg184 367 0 50.0000fF 
Lg184 367 368 57.0000pH
B184 367 368 10183 jj0 
Cgg184 368 0 50.0000fF
Vmeas184 368 369 0V

*Flux Biasing 
Idc185 0 50185 pwl(0 0uA 5ns 14.0680uA) 
Lflux185 50185 0 57.0000pH 
K185 Lg185 Lflux185 1

Cg185 369 0 50.0000fF 
Lg185 369 370 57.0000pH
B185 369 370 10184 jj0 
Cgg185 370 0 50.0000fF
Vmeas185 370 371 0V

*Flux Biasing 
Idc186 0 50186 pwl(0 0uA 5ns 14.0680uA) 
Lflux186 50186 0 57.0000pH 
K186 Lg186 Lflux186 1

Cg186 371 0 50.0000fF 
Lg186 371 372 57.0000pH
B186 371 372 10185 jj0 
Cgg186 372 0 50.0000fF
Vmeas186 372 373 0V

*Flux Biasing 
Idc187 0 50187 pwl(0 0uA 5ns 14.0680uA) 
Lflux187 50187 0 57.0000pH 
K187 Lg187 Lflux187 1

Cg187 373 0 50.0000fF 
Lg187 373 374 57.0000pH
B187 373 374 10186 jj0 
Cgg187 374 0 50.0000fF
Vmeas187 374 375 0V

*Flux Biasing 
Idc188 0 50188 pwl(0 0uA 5ns 14.0680uA) 
Lflux188 50188 0 57.0000pH 
K188 Lg188 Lflux188 1

Cg188 375 0 50.0000fF 
Lg188 375 376 57.0000pH
B188 375 376 10187 jj0 
Cgg188 376 0 50.0000fF
Vmeas188 376 377 0V

*Flux Biasing 
Idc189 0 50189 pwl(0 0uA 5ns 14.0680uA) 
Lflux189 50189 0 57.0000pH 
K189 Lg189 Lflux189 1

Cg189 377 0 50.0000fF 
Lg189 377 378 57.0000pH
B189 377 378 10188 jj0 
Cgg189 378 0 50.0000fF
Vmeas189 378 379 0V

*Flux Biasing 
Idc190 0 50190 pwl(0 0uA 5ns 14.0680uA) 
Lflux190 50190 0 57.0000pH 
K190 Lg190 Lflux190 1

Cg190 379 0 50.0000fF 
Lg190 379 380 57.0000pH
B190 379 380 10189 jj0 
Cgg190 380 0 50.0000fF
Vmeas190 380 381 0V

*Flux Biasing 
Idc191 0 50191 pwl(0 0uA 5ns 14.0680uA) 
Lflux191 50191 0 57.0000pH 
K191 Lg191 Lflux191 1

Cg191 381 0 50.0000fF 
Lg191 381 382 57.0000pH
B191 381 382 10190 jj0 
Cgg191 382 0 50.0000fF
Vmeas191 382 383 0V

*Flux Biasing 
Idc192 0 50192 pwl(0 0uA 5ns 14.0680uA) 
Lflux192 50192 0 57.0000pH 
K192 Lg192 Lflux192 1

Cg192 383 0 50.0000fF 
Lg192 383 384 57.0000pH
B192 383 384 10191 jj0 
Cgg192 384 0 50.0000fF
Vmeas192 384 385 0V

*Flux Biasing 
Idc193 0 50193 pwl(0 0uA 5ns 14.0680uA) 
Lflux193 50193 0 57.0000pH 
K193 Lg193 Lflux193 1

Cg193 385 0 50.0000fF 
Lg193 385 386 57.0000pH
B193 385 386 10192 jj0 
Cgg193 386 0 50.0000fF
Vmeas193 386 387 0V

*Flux Biasing 
Idc194 0 50194 pwl(0 0uA 5ns 14.0680uA) 
Lflux194 50194 0 57.0000pH 
K194 Lg194 Lflux194 1

Cg194 387 0 50.0000fF 
Lg194 387 388 57.0000pH
B194 387 388 10193 jj0 
Cgg194 388 0 50.0000fF
Vmeas194 388 389 0V

*Flux Biasing 
Idc195 0 50195 pwl(0 0uA 5ns 14.0680uA) 
Lflux195 50195 0 57.0000pH 
K195 Lg195 Lflux195 1

Cg195 389 0 50.0000fF 
Lg195 389 390 57.0000pH
B195 389 390 10194 jj0 
Cgg195 390 0 50.0000fF
Vmeas195 390 391 0V

*Flux Biasing 
Idc196 0 50196 pwl(0 0uA 5ns 14.0680uA) 
Lflux196 50196 0 57.0000pH 
K196 Lg196 Lflux196 1

Cg196 391 0 50.0000fF 
Lg196 391 392 57.0000pH
B196 391 392 10195 jj0 
Cgg196 392 0 50.0000fF
Vmeas196 392 393 0V

*Flux Biasing 
Idc197 0 50197 pwl(0 0uA 5ns 14.0680uA) 
Lflux197 50197 0 57.0000pH 
K197 Lg197 Lflux197 1

Cg197 393 0 50.0000fF 
Lg197 393 394 57.0000pH
B197 393 394 10196 jj0 
Cgg197 394 0 50.0000fF
Vmeas197 394 395 0V

*Flux Biasing 
Idc198 0 50198 pwl(0 0uA 5ns 14.0680uA) 
Lflux198 50198 0 57.0000pH 
K198 Lg198 Lflux198 1

Cg198 395 0 50.0000fF 
Lg198 395 396 57.0000pH
B198 395 396 10197 jj0 
Cgg198 396 0 50.0000fF
Vmeas198 396 397 0V

*Flux Biasing 
Idc199 0 50199 pwl(0 0uA 5ns 14.0680uA) 
Lflux199 50199 0 57.0000pH 
K199 Lg199 Lflux199 1

Cg199 397 0 50.0000fF 
Lg199 397 398 57.0000pH
B199 397 398 10198 jj0 
Cgg199 398 0 50.0000fF
Vmeas199 398 399 0V

*Flux Biasing 
Idc200 0 50200 pwl(0 0uA 5ns 14.0680uA) 
Lflux200 50200 0 57.0000pH 
K200 Lg200 Lflux200 1

Cg200 399 0 50.0000fF 
Lg200 399 400 57.0000pH
B200 399 400 10199 jj0 
Cgg200 400 0 50.0000fF
Vmeas200 400 401 0V

*Flux Biasing 
Idc201 0 50201 pwl(0 0uA 5ns 14.0680uA) 
Lflux201 50201 0 57.0000pH 
K201 Lg201 Lflux201 1

Cg201 401 0 50.0000fF 
Lg201 401 402 57.0000pH
B201 401 402 10200 jj0 
Cgg201 402 0 50.0000fF
Vmeas201 402 403 0V

*Flux Biasing 
Idc202 0 50202 pwl(0 0uA 5ns 14.0680uA) 
Lflux202 50202 0 57.0000pH 
K202 Lg202 Lflux202 1

Cg202 403 0 50.0000fF 
Lg202 403 404 57.0000pH
B202 403 404 10201 jj0 
Cgg202 404 0 50.0000fF
Vmeas202 404 405 0V

*Flux Biasing 
Idc203 0 50203 pwl(0 0uA 5ns 14.0680uA) 
Lflux203 50203 0 57.0000pH 
K203 Lg203 Lflux203 1

Cg203 405 0 50.0000fF 
Lg203 405 406 57.0000pH
B203 405 406 10202 jj0 
Cgg203 406 0 50.0000fF
Vmeas203 406 407 0V

*Flux Biasing 
Idc204 0 50204 pwl(0 0uA 5ns 14.0680uA) 
Lflux204 50204 0 57.0000pH 
K204 Lg204 Lflux204 1

Cg204 407 0 50.0000fF 
Lg204 407 408 57.0000pH
B204 407 408 10203 jj0 
Cgg204 408 0 50.0000fF
Vmeas204 408 409 0V

*Flux Biasing 
Idc205 0 50205 pwl(0 0uA 5ns 14.0680uA) 
Lflux205 50205 0 57.0000pH 
K205 Lg205 Lflux205 1

Cg205 409 0 50.0000fF 
Lg205 409 410 57.0000pH
B205 409 410 10204 jj0 
Cgg205 410 0 50.0000fF
Vmeas205 410 411 0V

*Flux Biasing 
Idc206 0 50206 pwl(0 0uA 5ns 14.0680uA) 
Lflux206 50206 0 57.0000pH 
K206 Lg206 Lflux206 1

Cg206 411 0 50.0000fF 
Lg206 411 412 57.0000pH
B206 411 412 10205 jj0 
Cgg206 412 0 50.0000fF
Vmeas206 412 413 0V

*Flux Biasing 
Idc207 0 50207 pwl(0 0uA 5ns 14.0680uA) 
Lflux207 50207 0 57.0000pH 
K207 Lg207 Lflux207 1

Cg207 413 0 50.0000fF 
Lg207 413 414 57.0000pH
B207 413 414 10206 jj0 
Cgg207 414 0 50.0000fF
Vmeas207 414 415 0V

*Flux Biasing 
Idc208 0 50208 pwl(0 0uA 5ns 14.0680uA) 
Lflux208 50208 0 57.0000pH 
K208 Lg208 Lflux208 1

Cg208 415 0 50.0000fF 
Lg208 415 416 57.0000pH
B208 415 416 10207 jj0 
Cgg208 416 0 50.0000fF
Vmeas208 416 417 0V

*Flux Biasing 
Idc209 0 50209 pwl(0 0uA 5ns 14.0680uA) 
Lflux209 50209 0 57.0000pH 
K209 Lg209 Lflux209 1

Cg209 417 0 50.0000fF 
Lg209 417 418 57.0000pH
B209 417 418 10208 jj0 
Cgg209 418 0 50.0000fF
Vmeas209 418 419 0V

*Flux Biasing 
Idc210 0 50210 pwl(0 0uA 5ns 14.0680uA) 
Lflux210 50210 0 57.0000pH 
K210 Lg210 Lflux210 1

Cg210 419 0 50.0000fF 
Lg210 419 420 57.0000pH
B210 419 420 10209 jj0 
Cgg210 420 0 50.0000fF
Vmeas210 420 421 0V

*Flux Biasing 
Idc211 0 50211 pwl(0 0uA 5ns 14.0680uA) 
Lflux211 50211 0 57.0000pH 
K211 Lg211 Lflux211 1

Cg211 421 0 50.0000fF 
Lg211 421 422 57.0000pH
B211 421 422 10210 jj0 
Cgg211 422 0 50.0000fF
Vmeas211 422 423 0V

*Flux Biasing 
Idc212 0 50212 pwl(0 0uA 5ns 14.0680uA) 
Lflux212 50212 0 57.0000pH 
K212 Lg212 Lflux212 1

Cg212 423 0 50.0000fF 
Lg212 423 424 57.0000pH
B212 423 424 10211 jj0 
Cgg212 424 0 50.0000fF
Vmeas212 424 425 0V

*Flux Biasing 
Idc213 0 50213 pwl(0 0uA 5ns 14.0680uA) 
Lflux213 50213 0 57.0000pH 
K213 Lg213 Lflux213 1

Cg213 425 0 50.0000fF 
Lg213 425 426 57.0000pH
B213 425 426 10212 jj0 
Cgg213 426 0 50.0000fF
Vmeas213 426 427 0V

*Flux Biasing 
Idc214 0 50214 pwl(0 0uA 5ns 14.0680uA) 
Lflux214 50214 0 57.0000pH 
K214 Lg214 Lflux214 1

Cg214 427 0 50.0000fF 
Lg214 427 428 57.0000pH
B214 427 428 10213 jj0 
Cgg214 428 0 50.0000fF
Vmeas214 428 429 0V

*Flux Biasing 
Idc215 0 50215 pwl(0 0uA 5ns 14.0680uA) 
Lflux215 50215 0 57.0000pH 
K215 Lg215 Lflux215 1

Cg215 429 0 50.0000fF 
Lg215 429 430 57.0000pH
B215 429 430 10214 jj0 
Cgg215 430 0 50.0000fF
Vmeas215 430 431 0V

*Flux Biasing 
Idc216 0 50216 pwl(0 0uA 5ns 14.0680uA) 
Lflux216 50216 0 57.0000pH 
K216 Lg216 Lflux216 1

Cg216 431 0 50.0000fF 
Lg216 431 432 57.0000pH
B216 431 432 10215 jj0 
Cgg216 432 0 50.0000fF
Vmeas216 432 433 0V

*Flux Biasing 
Idc217 0 50217 pwl(0 0uA 5ns 14.0680uA) 
Lflux217 50217 0 57.0000pH 
K217 Lg217 Lflux217 1

Cg217 433 0 50.0000fF 
Lg217 433 434 57.0000pH
B217 433 434 10216 jj0 
Cgg217 434 0 50.0000fF
Vmeas217 434 435 0V

*Flux Biasing 
Idc218 0 50218 pwl(0 0uA 5ns 14.0680uA) 
Lflux218 50218 0 57.0000pH 
K218 Lg218 Lflux218 1

Cg218 435 0 50.0000fF 
Lg218 435 436 57.0000pH
B218 435 436 10217 jj0 
Cgg218 436 0 50.0000fF
Vmeas218 436 437 0V

*Flux Biasing 
Idc219 0 50219 pwl(0 0uA 5ns 14.0680uA) 
Lflux219 50219 0 57.0000pH 
K219 Lg219 Lflux219 1

Cg219 437 0 50.0000fF 
Lg219 437 438 57.0000pH
B219 437 438 10218 jj0 
Cgg219 438 0 50.0000fF
Vmeas219 438 439 0V

*Flux Biasing 
Idc220 0 50220 pwl(0 0uA 5ns 14.0680uA) 
Lflux220 50220 0 57.0000pH 
K220 Lg220 Lflux220 1

Cg220 439 0 50.0000fF 
Lg220 439 440 57.0000pH
B220 439 440 10219 jj0 
Cgg220 440 0 50.0000fF
Vmeas220 440 441 0V

*Flux Biasing 
Idc221 0 50221 pwl(0 0uA 5ns 14.0680uA) 
Lflux221 50221 0 57.0000pH 
K221 Lg221 Lflux221 1

Cg221 441 0 50.0000fF 
Lg221 441 442 57.0000pH
B221 441 442 10220 jj0 
Cgg221 442 0 50.0000fF
Vmeas221 442 443 0V

*Flux Biasing 
Idc222 0 50222 pwl(0 0uA 5ns 14.0680uA) 
Lflux222 50222 0 57.0000pH 
K222 Lg222 Lflux222 1

Cg222 443 0 50.0000fF 
Lg222 443 444 57.0000pH
B222 443 444 10221 jj0 
Cgg222 444 0 50.0000fF
Vmeas222 444 445 0V

*Flux Biasing 
Idc223 0 50223 pwl(0 0uA 5ns 14.0680uA) 
Lflux223 50223 0 57.0000pH 
K223 Lg223 Lflux223 1

Cg223 445 0 50.0000fF 
Lg223 445 446 57.0000pH
B223 445 446 10222 jj0 
Cgg223 446 0 50.0000fF
Vmeas223 446 447 0V

*Flux Biasing 
Idc224 0 50224 pwl(0 0uA 5ns 14.0680uA) 
Lflux224 50224 0 57.0000pH 
K224 Lg224 Lflux224 1

Cg224 447 0 50.0000fF 
Lg224 447 448 57.0000pH
B224 447 448 10223 jj0 
Cgg224 448 0 50.0000fF
Vmeas224 448 449 0V

*Flux Biasing 
Idc225 0 50225 pwl(0 0uA 5ns 14.0680uA) 
Lflux225 50225 0 57.0000pH 
K225 Lg225 Lflux225 1

Cg225 449 0 50.0000fF 
Lg225 449 450 57.0000pH
B225 449 450 10224 jj0 
Cgg225 450 0 50.0000fF
Vmeas225 450 451 0V

*Flux Biasing 
Idc226 0 50226 pwl(0 0uA 5ns 14.0680uA) 
Lflux226 50226 0 57.0000pH 
K226 Lg226 Lflux226 1

Cg226 451 0 50.0000fF 
Lg226 451 452 57.0000pH
B226 451 452 10225 jj0 
Cgg226 452 0 50.0000fF
Vmeas226 452 453 0V

*Flux Biasing 
Idc227 0 50227 pwl(0 0uA 5ns 14.0680uA) 
Lflux227 50227 0 57.0000pH 
K227 Lg227 Lflux227 1

Cg227 453 0 50.0000fF 
Lg227 453 454 57.0000pH
B227 453 454 10226 jj0 
Cgg227 454 0 50.0000fF
Vmeas227 454 455 0V

*Flux Biasing 
Idc228 0 50228 pwl(0 0uA 5ns 14.0680uA) 
Lflux228 50228 0 57.0000pH 
K228 Lg228 Lflux228 1

Cg228 455 0 50.0000fF 
Lg228 455 456 57.0000pH
B228 455 456 10227 jj0 
Cgg228 456 0 50.0000fF
Vmeas228 456 457 0V

*Flux Biasing 
Idc229 0 50229 pwl(0 0uA 5ns 14.0680uA) 
Lflux229 50229 0 57.0000pH 
K229 Lg229 Lflux229 1

Cg229 457 0 50.0000fF 
Lg229 457 458 57.0000pH
B229 457 458 10228 jj0 
Cgg229 458 0 50.0000fF
Vmeas229 458 459 0V

*Flux Biasing 
Idc230 0 50230 pwl(0 0uA 5ns 14.0680uA) 
Lflux230 50230 0 57.0000pH 
K230 Lg230 Lflux230 1

Cg230 459 0 50.0000fF 
Lg230 459 460 57.0000pH
B230 459 460 10229 jj0 
Cgg230 460 0 50.0000fF
Vmeas230 460 461 0V

*Flux Biasing 
Idc231 0 50231 pwl(0 0uA 5ns 14.0680uA) 
Lflux231 50231 0 57.0000pH 
K231 Lg231 Lflux231 1

Cg231 461 0 50.0000fF 
Lg231 461 462 57.0000pH
B231 461 462 10230 jj0 
Cgg231 462 0 50.0000fF
Vmeas231 462 463 0V

*Flux Biasing 
Idc232 0 50232 pwl(0 0uA 5ns 14.0680uA) 
Lflux232 50232 0 57.0000pH 
K232 Lg232 Lflux232 1

Cg232 463 0 50.0000fF 
Lg232 463 464 57.0000pH
B232 463 464 10231 jj0 
Cgg232 464 0 50.0000fF
Vmeas232 464 465 0V

*Flux Biasing 
Idc233 0 50233 pwl(0 0uA 5ns 14.0680uA) 
Lflux233 50233 0 57.0000pH 
K233 Lg233 Lflux233 1

Cg233 465 0 50.0000fF 
Lg233 465 466 57.0000pH
B233 465 466 10232 jj0 
Cgg233 466 0 50.0000fF
Vmeas233 466 467 0V

*Flux Biasing 
Idc234 0 50234 pwl(0 0uA 5ns 14.0680uA) 
Lflux234 50234 0 57.0000pH 
K234 Lg234 Lflux234 1

Cg234 467 0 50.0000fF 
Lg234 467 468 57.0000pH
B234 467 468 10233 jj0 
Cgg234 468 0 50.0000fF
Vmeas234 468 469 0V

*Flux Biasing 
Idc235 0 50235 pwl(0 0uA 5ns 14.0680uA) 
Lflux235 50235 0 57.0000pH 
K235 Lg235 Lflux235 1

Cg235 469 0 50.0000fF 
Lg235 469 470 57.0000pH
B235 469 470 10234 jj0 
Cgg235 470 0 50.0000fF
Vmeas235 470 471 0V

*Flux Biasing 
Idc236 0 50236 pwl(0 0uA 5ns 14.0680uA) 
Lflux236 50236 0 57.0000pH 
K236 Lg236 Lflux236 1

Cg236 471 0 50.0000fF 
Lg236 471 472 57.0000pH
B236 471 472 10235 jj0 
Cgg236 472 0 50.0000fF
Vmeas236 472 473 0V

*Flux Biasing 
Idc237 0 50237 pwl(0 0uA 5ns 14.0680uA) 
Lflux237 50237 0 57.0000pH 
K237 Lg237 Lflux237 1

Cg237 473 0 50.0000fF 
Lg237 473 474 57.0000pH
B237 473 474 10236 jj0 
Cgg237 474 0 50.0000fF
Vmeas237 474 475 0V

*Flux Biasing 
Idc238 0 50238 pwl(0 0uA 5ns 14.0680uA) 
Lflux238 50238 0 57.0000pH 
K238 Lg238 Lflux238 1

Cg238 475 0 50.0000fF 
Lg238 475 476 57.0000pH
B238 475 476 10237 jj0 
Cgg238 476 0 50.0000fF
Vmeas238 476 477 0V

*Flux Biasing 
Idc239 0 50239 pwl(0 0uA 5ns 14.0680uA) 
Lflux239 50239 0 57.0000pH 
K239 Lg239 Lflux239 1

Cg239 477 0 50.0000fF 
Lg239 477 478 57.0000pH
B239 477 478 10238 jj0 
Cgg239 478 0 50.0000fF
Vmeas239 478 479 0V

*Flux Biasing 
Idc240 0 50240 pwl(0 0uA 5ns 14.0680uA) 
Lflux240 50240 0 57.0000pH 
K240 Lg240 Lflux240 1

Cg240 479 0 50.0000fF 
Lg240 479 480 57.0000pH
B240 479 480 10239 jj0 
Cgg240 480 0 50.0000fF
Vmeas240 480 481 0V

*Flux Biasing 
Idc241 0 50241 pwl(0 0uA 5ns 14.0680uA) 
Lflux241 50241 0 57.0000pH 
K241 Lg241 Lflux241 1

Cg241 481 0 50.0000fF 
Lg241 481 482 57.0000pH
B241 481 482 10240 jj0 
Cgg241 482 0 50.0000fF
Vmeas241 482 483 0V

*Flux Biasing 
Idc242 0 50242 pwl(0 0uA 5ns 14.0680uA) 
Lflux242 50242 0 57.0000pH 
K242 Lg242 Lflux242 1

Cg242 483 0 50.0000fF 
Lg242 483 484 57.0000pH
B242 483 484 10241 jj0 
Cgg242 484 0 50.0000fF
Vmeas242 484 485 0V

*Flux Biasing 
Idc243 0 50243 pwl(0 0uA 5ns 14.0680uA) 
Lflux243 50243 0 57.0000pH 
K243 Lg243 Lflux243 1

Cg243 485 0 50.0000fF 
Lg243 485 486 57.0000pH
B243 485 486 10242 jj0 
Cgg243 486 0 50.0000fF
Vmeas243 486 487 0V

*Flux Biasing 
Idc244 0 50244 pwl(0 0uA 5ns 14.0680uA) 
Lflux244 50244 0 57.0000pH 
K244 Lg244 Lflux244 1

Cg244 487 0 50.0000fF 
Lg244 487 488 57.0000pH
B244 487 488 10243 jj0 
Cgg244 488 0 50.0000fF
Vmeas244 488 489 0V

*Flux Biasing 
Idc245 0 50245 pwl(0 0uA 5ns 14.0680uA) 
Lflux245 50245 0 57.0000pH 
K245 Lg245 Lflux245 1

Cg245 489 0 50.0000fF 
Lg245 489 490 57.0000pH
B245 489 490 10244 jj0 
Cgg245 490 0 50.0000fF
Vmeas245 490 491 0V

*Flux Biasing 
Idc246 0 50246 pwl(0 0uA 5ns 14.0680uA) 
Lflux246 50246 0 57.0000pH 
K246 Lg246 Lflux246 1

Cg246 491 0 50.0000fF 
Lg246 491 492 57.0000pH
B246 491 492 10245 jj0 
Cgg246 492 0 50.0000fF
Vmeas246 492 493 0V

*Flux Biasing 
Idc247 0 50247 pwl(0 0uA 5ns 14.0680uA) 
Lflux247 50247 0 57.0000pH 
K247 Lg247 Lflux247 1

Cg247 493 0 50.0000fF 
Lg247 493 494 57.0000pH
B247 493 494 10246 jj0 
Cgg247 494 0 50.0000fF
Vmeas247 494 495 0V

*Flux Biasing 
Idc248 0 50248 pwl(0 0uA 5ns 14.0680uA) 
Lflux248 50248 0 57.0000pH 
K248 Lg248 Lflux248 1

Cg248 495 0 50.0000fF 
Lg248 495 496 57.0000pH
B248 495 496 10247 jj0 
Cgg248 496 0 50.0000fF
Vmeas248 496 497 0V

*Flux Biasing 
Idc249 0 50249 pwl(0 0uA 5ns 14.0680uA) 
Lflux249 50249 0 57.0000pH 
K249 Lg249 Lflux249 1

Cg249 497 0 50.0000fF 
Lg249 497 498 57.0000pH
B249 497 498 10248 jj0 
Cgg249 498 0 50.0000fF
Vmeas249 498 499 0V

*Flux Biasing 
Idc250 0 50250 pwl(0 0uA 5ns 14.0680uA) 
Lflux250 50250 0 57.0000pH 
K250 Lg250 Lflux250 1

Cg250 499 0 50.0000fF 
Lg250 499 500 57.0000pH
B250 499 500 10249 jj0 
Cgg250 500 0 50.0000fF
Vmeas250 500 501 0V

*Flux Biasing 
Idc251 0 50251 pwl(0 0uA 5ns 14.0680uA) 
Lflux251 50251 0 57.0000pH 
K251 Lg251 Lflux251 1

Cg251 501 0 50.0000fF 
Lg251 501 502 57.0000pH
B251 501 502 10250 jj0 
Cgg251 502 0 50.0000fF
Vmeas251 502 503 0V

*Flux Biasing 
Idc252 0 50252 pwl(0 0uA 5ns 14.0680uA) 
Lflux252 50252 0 57.0000pH 
K252 Lg252 Lflux252 1

Cg252 503 0 50.0000fF 
Lg252 503 504 57.0000pH
B252 503 504 10251 jj0 
Cgg252 504 0 50.0000fF
Vmeas252 504 505 0V

*Flux Biasing 
Idc253 0 50253 pwl(0 0uA 5ns 14.0680uA) 
Lflux253 50253 0 57.0000pH 
K253 Lg253 Lflux253 1

Cg253 505 0 50.0000fF 
Lg253 505 506 57.0000pH
B253 505 506 10252 jj0 
Cgg253 506 0 50.0000fF
Vmeas253 506 507 0V

*Flux Biasing 
Idc254 0 50254 pwl(0 0uA 5ns 14.0680uA) 
Lflux254 50254 0 57.0000pH 
K254 Lg254 Lflux254 1

Cg254 507 0 50.0000fF 
Lg254 507 508 57.0000pH
B254 507 508 10253 jj0 
Cgg254 508 0 50.0000fF
Vmeas254 508 509 0V

*Flux Biasing 
Idc255 0 50255 pwl(0 0uA 5ns 14.0680uA) 
Lflux255 50255 0 57.0000pH 
K255 Lg255 Lflux255 1

Cg255 509 0 50.0000fF 
Lg255 509 510 57.0000pH
B255 509 510 10254 jj0 
Cgg255 510 0 50.0000fF
Vmeas255 510 511 0V

*Flux Biasing 
Idc256 0 50256 pwl(0 0uA 5ns 14.0680uA) 
Lflux256 50256 0 57.0000pH 
K256 Lg256 Lflux256 1

Cg256 511 0 50.0000fF 
Lg256 511 512 57.0000pH
B256 511 512 10255 jj0 
Cgg256 512 0 50.0000fF
Vmeas256 512 513 0V

*Flux Biasing 
Idc257 0 50257 pwl(0 0uA 5ns 14.0680uA) 
Lflux257 50257 0 57.0000pH 
K257 Lg257 Lflux257 1

Cg257 513 0 50.0000fF 
Lg257 513 514 57.0000pH
B257 513 514 10256 jj0 
Cgg257 514 0 50.0000fF
Vmeas257 514 515 0V

*Flux Biasing 
Idc258 0 50258 pwl(0 0uA 5ns 14.0680uA) 
Lflux258 50258 0 57.0000pH 
K258 Lg258 Lflux258 1

Cg258 515 0 50.0000fF 
Lg258 515 516 57.0000pH
B258 515 516 10257 jj0 
Cgg258 516 0 50.0000fF
Vmeas258 516 517 0V

*Flux Biasing 
Idc259 0 50259 pwl(0 0uA 5ns 14.0680uA) 
Lflux259 50259 0 57.0000pH 
K259 Lg259 Lflux259 1

Cg259 517 0 50.0000fF 
Lg259 517 518 57.0000pH
B259 517 518 10258 jj0 
Cgg259 518 0 50.0000fF
Vmeas259 518 519 0V

*Flux Biasing 
Idc260 0 50260 pwl(0 0uA 5ns 14.0680uA) 
Lflux260 50260 0 57.0000pH 
K260 Lg260 Lflux260 1

Cg260 519 0 50.0000fF 
Lg260 519 520 57.0000pH
B260 519 520 10259 jj0 
Cgg260 520 0 50.0000fF
Vmeas260 520 521 0V

*Flux Biasing 
Idc261 0 50261 pwl(0 0uA 5ns 14.0680uA) 
Lflux261 50261 0 57.0000pH 
K261 Lg261 Lflux261 1

Cg261 521 0 50.0000fF 
Lg261 521 522 57.0000pH
B261 521 522 10260 jj0 
Cgg261 522 0 50.0000fF
Vmeas261 522 523 0V

*Flux Biasing 
Idc262 0 50262 pwl(0 0uA 5ns 14.0680uA) 
Lflux262 50262 0 57.0000pH 
K262 Lg262 Lflux262 1

Cg262 523 0 50.0000fF 
Lg262 523 524 57.0000pH
B262 523 524 10261 jj0 
Cgg262 524 0 50.0000fF
Vmeas262 524 525 0V

*Flux Biasing 
Idc263 0 50263 pwl(0 0uA 5ns 14.0680uA) 
Lflux263 50263 0 57.0000pH 
K263 Lg263 Lflux263 1

Cg263 525 0 50.0000fF 
Lg263 525 526 57.0000pH
B263 525 526 10262 jj0 
Cgg263 526 0 50.0000fF
Vmeas263 526 527 0V

*Flux Biasing 
Idc264 0 50264 pwl(0 0uA 5ns 14.0680uA) 
Lflux264 50264 0 57.0000pH 
K264 Lg264 Lflux264 1

Cg264 527 0 50.0000fF 
Lg264 527 528 57.0000pH
B264 527 528 10263 jj0 
Cgg264 528 0 50.0000fF
Vmeas264 528 529 0V

*Flux Biasing 
Idc265 0 50265 pwl(0 0uA 5ns 14.0680uA) 
Lflux265 50265 0 57.0000pH 
K265 Lg265 Lflux265 1

Cg265 529 0 50.0000fF 
Lg265 529 530 57.0000pH
B265 529 530 10264 jj0 
Cgg265 530 0 50.0000fF
Vmeas265 530 531 0V

*Flux Biasing 
Idc266 0 50266 pwl(0 0uA 5ns 14.0680uA) 
Lflux266 50266 0 57.0000pH 
K266 Lg266 Lflux266 1

Cg266 531 0 50.0000fF 
Lg266 531 532 57.0000pH
B266 531 532 10265 jj0 
Cgg266 532 0 50.0000fF
Vmeas266 532 533 0V

*Flux Biasing 
Idc267 0 50267 pwl(0 0uA 5ns 14.0680uA) 
Lflux267 50267 0 57.0000pH 
K267 Lg267 Lflux267 1

Cg267 533 0 50.0000fF 
Lg267 533 534 57.0000pH
B267 533 534 10266 jj0 
Cgg267 534 0 50.0000fF
Vmeas267 534 535 0V

*Flux Biasing 
Idc268 0 50268 pwl(0 0uA 5ns 14.0680uA) 
Lflux268 50268 0 57.0000pH 
K268 Lg268 Lflux268 1

Cg268 535 0 50.0000fF 
Lg268 535 536 57.0000pH
B268 535 536 10267 jj0 
Cgg268 536 0 50.0000fF
Vmeas268 536 537 0V

*Flux Biasing 
Idc269 0 50269 pwl(0 0uA 5ns 14.0680uA) 
Lflux269 50269 0 57.0000pH 
K269 Lg269 Lflux269 1

Cg269 537 0 50.0000fF 
Lg269 537 538 57.0000pH
B269 537 538 10268 jj0 
Cgg269 538 0 50.0000fF
Vmeas269 538 539 0V

*Flux Biasing 
Idc270 0 50270 pwl(0 0uA 5ns 14.0680uA) 
Lflux270 50270 0 57.0000pH 
K270 Lg270 Lflux270 1

Cg270 539 0 50.0000fF 
Lg270 539 540 57.0000pH
B270 539 540 10269 jj0 
Cgg270 540 0 50.0000fF
Vmeas270 540 541 0V

*Flux Biasing 
Idc271 0 50271 pwl(0 0uA 5ns 14.0680uA) 
Lflux271 50271 0 57.0000pH 
K271 Lg271 Lflux271 1

Cg271 541 0 50.0000fF 
Lg271 541 542 57.0000pH
B271 541 542 10270 jj0 
Cgg271 542 0 50.0000fF
Vmeas271 542 543 0V

*Flux Biasing 
Idc272 0 50272 pwl(0 0uA 5ns 14.0680uA) 
Lflux272 50272 0 57.0000pH 
K272 Lg272 Lflux272 1

Cg272 543 0 50.0000fF 
Lg272 543 544 57.0000pH
B272 543 544 10271 jj0 
Cgg272 544 0 50.0000fF
Vmeas272 544 545 0V

*Flux Biasing 
Idc273 0 50273 pwl(0 0uA 5ns 14.0680uA) 
Lflux273 50273 0 57.0000pH 
K273 Lg273 Lflux273 1

Cg273 545 0 50.0000fF 
Lg273 545 546 57.0000pH
B273 545 546 10272 jj0 
Cgg273 546 0 50.0000fF
Vmeas273 546 547 0V

*Flux Biasing 
Idc274 0 50274 pwl(0 0uA 5ns 14.0680uA) 
Lflux274 50274 0 57.0000pH 
K274 Lg274 Lflux274 1

Cg274 547 0 50.0000fF 
Lg274 547 548 57.0000pH
B274 547 548 10273 jj0 
Cgg274 548 0 50.0000fF
Vmeas274 548 549 0V

*Flux Biasing 
Idc275 0 50275 pwl(0 0uA 5ns 14.0680uA) 
Lflux275 50275 0 57.0000pH 
K275 Lg275 Lflux275 1

Cg275 549 0 50.0000fF 
Lg275 549 550 57.0000pH
B275 549 550 10274 jj0 
Cgg275 550 0 50.0000fF
Vmeas275 550 551 0V

*Flux Biasing 
Idc276 0 50276 pwl(0 0uA 5ns 14.0680uA) 
Lflux276 50276 0 57.0000pH 
K276 Lg276 Lflux276 1

Cg276 551 0 50.0000fF 
Lg276 551 552 57.0000pH
B276 551 552 10275 jj0 
Cgg276 552 0 50.0000fF
Vmeas276 552 553 0V

*Flux Biasing 
Idc277 0 50277 pwl(0 0uA 5ns 14.0680uA) 
Lflux277 50277 0 57.0000pH 
K277 Lg277 Lflux277 1

Cg277 553 0 50.0000fF 
Lg277 553 554 57.0000pH
B277 553 554 10276 jj0 
Cgg277 554 0 50.0000fF
Vmeas277 554 555 0V

*Flux Biasing 
Idc278 0 50278 pwl(0 0uA 5ns 14.0680uA) 
Lflux278 50278 0 57.0000pH 
K278 Lg278 Lflux278 1

Cg278 555 0 50.0000fF 
Lg278 555 556 57.0000pH
B278 555 556 10277 jj0 
Cgg278 556 0 50.0000fF
Vmeas278 556 557 0V

*Flux Biasing 
Idc279 0 50279 pwl(0 0uA 5ns 14.0680uA) 
Lflux279 50279 0 57.0000pH 
K279 Lg279 Lflux279 1

Cg279 557 0 50.0000fF 
Lg279 557 558 57.0000pH
B279 557 558 10278 jj0 
Cgg279 558 0 50.0000fF
Vmeas279 558 559 0V

*Flux Biasing 
Idc280 0 50280 pwl(0 0uA 5ns 14.0680uA) 
Lflux280 50280 0 57.0000pH 
K280 Lg280 Lflux280 1

Cg280 559 0 50.0000fF 
Lg280 559 560 57.0000pH
B280 559 560 10279 jj0 
Cgg280 560 0 50.0000fF
Vmeas280 560 561 0V

*Flux Biasing 
Idc281 0 50281 pwl(0 0uA 5ns 14.0680uA) 
Lflux281 50281 0 57.0000pH 
K281 Lg281 Lflux281 1

Cg281 561 0 50.0000fF 
Lg281 561 562 57.0000pH
B281 561 562 10280 jj0 
Cgg281 562 0 50.0000fF
Vmeas281 562 563 0V

*Flux Biasing 
Idc282 0 50282 pwl(0 0uA 5ns 14.0680uA) 
Lflux282 50282 0 57.0000pH 
K282 Lg282 Lflux282 1

Cg282 563 0 50.0000fF 
Lg282 563 564 57.0000pH
B282 563 564 10281 jj0 
Cgg282 564 0 50.0000fF
Vmeas282 564 565 0V

*Flux Biasing 
Idc283 0 50283 pwl(0 0uA 5ns 14.0680uA) 
Lflux283 50283 0 57.0000pH 
K283 Lg283 Lflux283 1

Cg283 565 0 50.0000fF 
Lg283 565 566 57.0000pH
B283 565 566 10282 jj0 
Cgg283 566 0 50.0000fF
Vmeas283 566 567 0V

*Flux Biasing 
Idc284 0 50284 pwl(0 0uA 5ns 14.0680uA) 
Lflux284 50284 0 57.0000pH 
K284 Lg284 Lflux284 1

Cg284 567 0 50.0000fF 
Lg284 567 568 57.0000pH
B284 567 568 10283 jj0 
Cgg284 568 0 50.0000fF
Vmeas284 568 569 0V

*Flux Biasing 
Idc285 0 50285 pwl(0 0uA 5ns 14.0680uA) 
Lflux285 50285 0 57.0000pH 
K285 Lg285 Lflux285 1

Cg285 569 0 50.0000fF 
Lg285 569 570 57.0000pH
B285 569 570 10284 jj0 
Cgg285 570 0 50.0000fF
Vmeas285 570 571 0V

*Flux Biasing 
Idc286 0 50286 pwl(0 0uA 5ns 14.0680uA) 
Lflux286 50286 0 57.0000pH 
K286 Lg286 Lflux286 1

Cg286 571 0 50.0000fF 
Lg286 571 572 57.0000pH
B286 571 572 10285 jj0 
Cgg286 572 0 50.0000fF
Vmeas286 572 573 0V

*Flux Biasing 
Idc287 0 50287 pwl(0 0uA 5ns 14.0680uA) 
Lflux287 50287 0 57.0000pH 
K287 Lg287 Lflux287 1

Cg287 573 0 50.0000fF 
Lg287 573 574 57.0000pH
B287 573 574 10286 jj0 
Cgg287 574 0 50.0000fF
Vmeas287 574 575 0V

*Flux Biasing 
Idc288 0 50288 pwl(0 0uA 5ns 14.0680uA) 
Lflux288 50288 0 57.0000pH 
K288 Lg288 Lflux288 1

Cg288 575 0 50.0000fF 
Lg288 575 576 57.0000pH
B288 575 576 10287 jj0 
Cgg288 576 0 50.0000fF
Vmeas288 576 577 0V

*Flux Biasing 
Idc289 0 50289 pwl(0 0uA 5ns 14.0680uA) 
Lflux289 50289 0 57.0000pH 
K289 Lg289 Lflux289 1

Cg289 577 0 50.0000fF 
Lg289 577 578 57.0000pH
B289 577 578 10288 jj0 
Cgg289 578 0 50.0000fF
Vmeas289 578 579 0V

*Flux Biasing 
Idc290 0 50290 pwl(0 0uA 5ns 14.0680uA) 
Lflux290 50290 0 57.0000pH 
K290 Lg290 Lflux290 1

Cg290 579 0 50.0000fF 
Lg290 579 580 57.0000pH
B290 579 580 10289 jj0 
Cgg290 580 0 50.0000fF
Vmeas290 580 581 0V

*Flux Biasing 
Idc291 0 50291 pwl(0 0uA 5ns 14.0680uA) 
Lflux291 50291 0 57.0000pH 
K291 Lg291 Lflux291 1

Cg291 581 0 50.0000fF 
Lg291 581 582 57.0000pH
B291 581 582 10290 jj0 
Cgg291 582 0 50.0000fF
Vmeas291 582 583 0V

*Flux Biasing 
Idc292 0 50292 pwl(0 0uA 5ns 14.0680uA) 
Lflux292 50292 0 57.0000pH 
K292 Lg292 Lflux292 1

Cg292 583 0 50.0000fF 
Lg292 583 584 57.0000pH
B292 583 584 10291 jj0 
Cgg292 584 0 50.0000fF
Vmeas292 584 585 0V

*Flux Biasing 
Idc293 0 50293 pwl(0 0uA 5ns 14.0680uA) 
Lflux293 50293 0 57.0000pH 
K293 Lg293 Lflux293 1

Cg293 585 0 50.0000fF 
Lg293 585 586 57.0000pH
B293 585 586 10292 jj0 
Cgg293 586 0 50.0000fF
Vmeas293 586 587 0V

*Flux Biasing 
Idc294 0 50294 pwl(0 0uA 5ns 14.0680uA) 
Lflux294 50294 0 57.0000pH 
K294 Lg294 Lflux294 1

Cg294 587 0 50.0000fF 
Lg294 587 588 57.0000pH
B294 587 588 10293 jj0 
Cgg294 588 0 50.0000fF
Vmeas294 588 589 0V

*Flux Biasing 
Idc295 0 50295 pwl(0 0uA 5ns 14.0680uA) 
Lflux295 50295 0 57.0000pH 
K295 Lg295 Lflux295 1

Cg295 589 0 50.0000fF 
Lg295 589 590 57.0000pH
B295 589 590 10294 jj0 
Cgg295 590 0 50.0000fF
Vmeas295 590 591 0V

*Flux Biasing 
Idc296 0 50296 pwl(0 0uA 5ns 14.0680uA) 
Lflux296 50296 0 57.0000pH 
K296 Lg296 Lflux296 1

Cg296 591 0 50.0000fF 
Lg296 591 592 57.0000pH
B296 591 592 10295 jj0 
Cgg296 592 0 50.0000fF
Vmeas296 592 593 0V

*Flux Biasing 
Idc297 0 50297 pwl(0 0uA 5ns 14.0680uA) 
Lflux297 50297 0 57.0000pH 
K297 Lg297 Lflux297 1

Cg297 593 0 50.0000fF 
Lg297 593 594 57.0000pH
B297 593 594 10296 jj0 
Cgg297 594 0 50.0000fF
Vmeas297 594 595 0V

*Flux Biasing 
Idc298 0 50298 pwl(0 0uA 5ns 14.0680uA) 
Lflux298 50298 0 57.0000pH 
K298 Lg298 Lflux298 1

Cg298 595 0 50.0000fF 
Lg298 595 596 57.0000pH
B298 595 596 10297 jj0 
Cgg298 596 0 50.0000fF
Vmeas298 596 597 0V

*Flux Biasing 
Idc299 0 50299 pwl(0 0uA 5ns 14.0680uA) 
Lflux299 50299 0 57.0000pH 
K299 Lg299 Lflux299 1

Cg299 597 0 50.0000fF 
Lg299 597 598 57.0000pH
B299 597 598 10298 jj0 
Cgg299 598 0 50.0000fF
Vmeas299 598 599 0V

*Flux Biasing 
Idc300 0 50300 pwl(0 0uA 5ns 14.0680uA) 
Lflux300 50300 0 57.0000pH 
K300 Lg300 Lflux300 1

Cg300 599 0 50.0000fF 
Lg300 599 600 57.0000pH
B300 599 600 10299 jj0 
Cgg300 600 0 50.0000fF
Vmeas300 600 601 0V

*Flux Biasing 
Idc301 0 50301 pwl(0 0uA 5ns 14.0680uA) 
Lflux301 50301 0 57.0000pH 
K301 Lg301 Lflux301 1

Cg301 601 0 50.0000fF 
Lg301 601 602 57.0000pH
B301 601 602 10300 jj0 
Cgg301 602 0 50.0000fF
Vmeas301 602 603 0V

*Flux Biasing 
Idc302 0 50302 pwl(0 0uA 5ns 14.0680uA) 
Lflux302 50302 0 57.0000pH 
K302 Lg302 Lflux302 1

Cg302 603 0 50.0000fF 
Lg302 603 604 57.0000pH
B302 603 604 10301 jj0 
Cgg302 604 0 50.0000fF
Vmeas302 604 605 0V

*Flux Biasing 
Idc303 0 50303 pwl(0 0uA 5ns 14.0680uA) 
Lflux303 50303 0 57.0000pH 
K303 Lg303 Lflux303 1

Cg303 605 0 50.0000fF 
Lg303 605 606 57.0000pH
B303 605 606 10302 jj0 
Cgg303 606 0 50.0000fF
Vmeas303 606 607 0V

*Flux Biasing 
Idc304 0 50304 pwl(0 0uA 5ns 14.0680uA) 
Lflux304 50304 0 57.0000pH 
K304 Lg304 Lflux304 1

Cg304 607 0 50.0000fF 
Lg304 607 608 57.0000pH
B304 607 608 10303 jj0 
Cgg304 608 0 50.0000fF
Vmeas304 608 609 0V

*Flux Biasing 
Idc305 0 50305 pwl(0 0uA 5ns 14.0680uA) 
Lflux305 50305 0 57.0000pH 
K305 Lg305 Lflux305 1

Cg305 609 0 50.0000fF 
Lg305 609 610 57.0000pH
B305 609 610 10304 jj0 
Cgg305 610 0 50.0000fF
Vmeas305 610 611 0V

*Flux Biasing 
Idc306 0 50306 pwl(0 0uA 5ns 14.0680uA) 
Lflux306 50306 0 57.0000pH 
K306 Lg306 Lflux306 1

Cg306 611 0 50.0000fF 
Lg306 611 612 57.0000pH
B306 611 612 10305 jj0 
Cgg306 612 0 50.0000fF
Vmeas306 612 613 0V

*Flux Biasing 
Idc307 0 50307 pwl(0 0uA 5ns 14.0680uA) 
Lflux307 50307 0 57.0000pH 
K307 Lg307 Lflux307 1

Cg307 613 0 50.0000fF 
Lg307 613 614 57.0000pH
B307 613 614 10306 jj0 
Cgg307 614 0 50.0000fF
Vmeas307 614 615 0V

*Flux Biasing 
Idc308 0 50308 pwl(0 0uA 5ns 14.0680uA) 
Lflux308 50308 0 57.0000pH 
K308 Lg308 Lflux308 1

Cg308 615 0 50.0000fF 
Lg308 615 616 57.0000pH
B308 615 616 10307 jj0 
Cgg308 616 0 50.0000fF
Vmeas308 616 617 0V

*Flux Biasing 
Idc309 0 50309 pwl(0 0uA 5ns 14.0680uA) 
Lflux309 50309 0 57.0000pH 
K309 Lg309 Lflux309 1

Cg309 617 0 50.0000fF 
Lg309 617 618 57.0000pH
B309 617 618 10308 jj0 
Cgg309 618 0 50.0000fF
Vmeas309 618 619 0V

*Flux Biasing 
Idc310 0 50310 pwl(0 0uA 5ns 14.0680uA) 
Lflux310 50310 0 57.0000pH 
K310 Lg310 Lflux310 1

Cg310 619 0 50.0000fF 
Lg310 619 620 57.0000pH
B310 619 620 10309 jj0 
Cgg310 620 0 50.0000fF
Vmeas310 620 621 0V

*Flux Biasing 
Idc311 0 50311 pwl(0 0uA 5ns 14.0680uA) 
Lflux311 50311 0 57.0000pH 
K311 Lg311 Lflux311 1

Cg311 621 0 50.0000fF 
Lg311 621 622 57.0000pH
B311 621 622 10310 jj0 
Cgg311 622 0 50.0000fF
Vmeas311 622 623 0V

*Flux Biasing 
Idc312 0 50312 pwl(0 0uA 5ns 14.0680uA) 
Lflux312 50312 0 57.0000pH 
K312 Lg312 Lflux312 1

Cg312 623 0 50.0000fF 
Lg312 623 624 57.0000pH
B312 623 624 10311 jj0 
Cgg312 624 0 50.0000fF
Vmeas312 624 625 0V

*Flux Biasing 
Idc313 0 50313 pwl(0 0uA 5ns 14.0680uA) 
Lflux313 50313 0 57.0000pH 
K313 Lg313 Lflux313 1

Cg313 625 0 50.0000fF 
Lg313 625 626 57.0000pH
B313 625 626 10312 jj0 
Cgg313 626 0 50.0000fF
Vmeas313 626 627 0V

*Flux Biasing 
Idc314 0 50314 pwl(0 0uA 5ns 14.0680uA) 
Lflux314 50314 0 57.0000pH 
K314 Lg314 Lflux314 1

Cg314 627 0 50.0000fF 
Lg314 627 628 57.0000pH
B314 627 628 10313 jj0 
Cgg314 628 0 50.0000fF
Vmeas314 628 629 0V

*Flux Biasing 
Idc315 0 50315 pwl(0 0uA 5ns 14.0680uA) 
Lflux315 50315 0 57.0000pH 
K315 Lg315 Lflux315 1

Cg315 629 0 50.0000fF 
Lg315 629 630 57.0000pH
B315 629 630 10314 jj0 
Cgg315 630 0 50.0000fF
Vmeas315 630 631 0V

*Flux Biasing 
Idc316 0 50316 pwl(0 0uA 5ns 14.0680uA) 
Lflux316 50316 0 57.0000pH 
K316 Lg316 Lflux316 1

Cg316 631 0 50.0000fF 
Lg316 631 632 57.0000pH
B316 631 632 10315 jj0 
Cgg316 632 0 50.0000fF
Vmeas316 632 633 0V

*Flux Biasing 
Idc317 0 50317 pwl(0 0uA 5ns 14.0680uA) 
Lflux317 50317 0 57.0000pH 
K317 Lg317 Lflux317 1

Cg317 633 0 50.0000fF 
Lg317 633 634 57.0000pH
B317 633 634 10316 jj0 
Cgg317 634 0 50.0000fF
Vmeas317 634 635 0V

*Flux Biasing 
Idc318 0 50318 pwl(0 0uA 5ns 14.0680uA) 
Lflux318 50318 0 57.0000pH 
K318 Lg318 Lflux318 1

Cg318 635 0 50.0000fF 
Lg318 635 636 57.0000pH
B318 635 636 10317 jj0 
Cgg318 636 0 50.0000fF
Vmeas318 636 637 0V

*Flux Biasing 
Idc319 0 50319 pwl(0 0uA 5ns 14.0680uA) 
Lflux319 50319 0 57.0000pH 
K319 Lg319 Lflux319 1

Cg319 637 0 50.0000fF 
Lg319 637 638 57.0000pH
B319 637 638 10318 jj0 
Cgg319 638 0 50.0000fF
Vmeas319 638 639 0V

*Flux Biasing 
Idc320 0 50320 pwl(0 0uA 5ns 14.0680uA) 
Lflux320 50320 0 57.0000pH 
K320 Lg320 Lflux320 1

Cg320 639 0 50.0000fF 
Lg320 639 640 57.0000pH
B320 639 640 10319 jj0 
Cgg320 640 0 50.0000fF
Vmeas320 640 641 0V

*Flux Biasing 
Idc321 0 50321 pwl(0 0uA 5ns 14.0680uA) 
Lflux321 50321 0 57.0000pH 
K321 Lg321 Lflux321 1

Cg321 641 0 50.0000fF 
Lg321 641 642 57.0000pH
B321 641 642 10320 jj0 
Cgg321 642 0 50.0000fF
Vmeas321 642 643 0V

*Flux Biasing 
Idc322 0 50322 pwl(0 0uA 5ns 14.0680uA) 
Lflux322 50322 0 57.0000pH 
K322 Lg322 Lflux322 1

Cg322 643 0 50.0000fF 
Lg322 643 644 57.0000pH
B322 643 644 10321 jj0 
Cgg322 644 0 50.0000fF
Vmeas322 644 645 0V

*Flux Biasing 
Idc323 0 50323 pwl(0 0uA 5ns 14.0680uA) 
Lflux323 50323 0 57.0000pH 
K323 Lg323 Lflux323 1

Cg323 645 0 50.0000fF 
Lg323 645 646 57.0000pH
B323 645 646 10322 jj0 
Cgg323 646 0 50.0000fF
Vmeas323 646 647 0V

*Flux Biasing 
Idc324 0 50324 pwl(0 0uA 5ns 14.0680uA) 
Lflux324 50324 0 57.0000pH 
K324 Lg324 Lflux324 1

Cg324 647 0 50.0000fF 
Lg324 647 648 57.0000pH
B324 647 648 10323 jj0 
Cgg324 648 0 50.0000fF
Vmeas324 648 649 0V

*Flux Biasing 
Idc325 0 50325 pwl(0 0uA 5ns 14.0680uA) 
Lflux325 50325 0 57.0000pH 
K325 Lg325 Lflux325 1

Cg325 649 0 50.0000fF 
Lg325 649 650 57.0000pH
B325 649 650 10324 jj0 
Cgg325 650 0 50.0000fF
Vmeas325 650 651 0V

*Flux Biasing 
Idc326 0 50326 pwl(0 0uA 5ns 14.0680uA) 
Lflux326 50326 0 57.0000pH 
K326 Lg326 Lflux326 1

Cg326 651 0 50.0000fF 
Lg326 651 652 57.0000pH
B326 651 652 10325 jj0 
Cgg326 652 0 50.0000fF
Vmeas326 652 653 0V

*Flux Biasing 
Idc327 0 50327 pwl(0 0uA 5ns 14.0680uA) 
Lflux327 50327 0 57.0000pH 
K327 Lg327 Lflux327 1

Cg327 653 0 50.0000fF 
Lg327 653 654 57.0000pH
B327 653 654 10326 jj0 
Cgg327 654 0 50.0000fF
Vmeas327 654 655 0V

*Flux Biasing 
Idc328 0 50328 pwl(0 0uA 5ns 14.0680uA) 
Lflux328 50328 0 57.0000pH 
K328 Lg328 Lflux328 1

Cg328 655 0 50.0000fF 
Lg328 655 656 57.0000pH
B328 655 656 10327 jj0 
Cgg328 656 0 50.0000fF
Vmeas328 656 657 0V

*Flux Biasing 
Idc329 0 50329 pwl(0 0uA 5ns 14.0680uA) 
Lflux329 50329 0 57.0000pH 
K329 Lg329 Lflux329 1

Cg329 657 0 50.0000fF 
Lg329 657 658 57.0000pH
B329 657 658 10328 jj0 
Cgg329 658 0 50.0000fF
Vmeas329 658 659 0V

*Flux Biasing 
Idc330 0 50330 pwl(0 0uA 5ns 14.0680uA) 
Lflux330 50330 0 57.0000pH 
K330 Lg330 Lflux330 1

Cg330 659 0 50.0000fF 
Lg330 659 660 57.0000pH
B330 659 660 10329 jj0 
Cgg330 660 0 50.0000fF
Vmeas330 660 661 0V

*Flux Biasing 
Idc331 0 50331 pwl(0 0uA 5ns 14.0680uA) 
Lflux331 50331 0 57.0000pH 
K331 Lg331 Lflux331 1

Cg331 661 0 50.0000fF 
Lg331 661 662 57.0000pH
B331 661 662 10330 jj0 
Cgg331 662 0 50.0000fF
Vmeas331 662 663 0V

*Flux Biasing 
Idc332 0 50332 pwl(0 0uA 5ns 14.0680uA) 
Lflux332 50332 0 57.0000pH 
K332 Lg332 Lflux332 1

Cg332 663 0 50.0000fF 
Lg332 663 664 57.0000pH
B332 663 664 10331 jj0 
Cgg332 664 0 50.0000fF
Vmeas332 664 665 0V

*Flux Biasing 
Idc333 0 50333 pwl(0 0uA 5ns 14.0680uA) 
Lflux333 50333 0 57.0000pH 
K333 Lg333 Lflux333 1

Cg333 665 0 50.0000fF 
Lg333 665 666 57.0000pH
B333 665 666 10332 jj0 
Cgg333 666 0 50.0000fF
Vmeas333 666 667 0V

*Flux Biasing 
Idc334 0 50334 pwl(0 0uA 5ns 14.0680uA) 
Lflux334 50334 0 57.0000pH 
K334 Lg334 Lflux334 1

Cg334 667 0 50.0000fF 
Lg334 667 668 57.0000pH
B334 667 668 10333 jj0 
Cgg334 668 0 50.0000fF
Vmeas334 668 669 0V

*Flux Biasing 
Idc335 0 50335 pwl(0 0uA 5ns 14.0680uA) 
Lflux335 50335 0 57.0000pH 
K335 Lg335 Lflux335 1

Cg335 669 0 50.0000fF 
Lg335 669 670 57.0000pH
B335 669 670 10334 jj0 
Cgg335 670 0 50.0000fF
Vmeas335 670 671 0V

*Flux Biasing 
Idc336 0 50336 pwl(0 0uA 5ns 14.0680uA) 
Lflux336 50336 0 57.0000pH 
K336 Lg336 Lflux336 1

Cg336 671 0 50.0000fF 
Lg336 671 672 57.0000pH
B336 671 672 10335 jj0 
Cgg336 672 0 50.0000fF
Vmeas336 672 673 0V

*Flux Biasing 
Idc337 0 50337 pwl(0 0uA 5ns 14.0680uA) 
Lflux337 50337 0 57.0000pH 
K337 Lg337 Lflux337 1

Cg337 673 0 50.0000fF 
Lg337 673 674 57.0000pH
B337 673 674 10336 jj0 
Cgg337 674 0 50.0000fF
Vmeas337 674 675 0V

*Flux Biasing 
Idc338 0 50338 pwl(0 0uA 5ns 14.0680uA) 
Lflux338 50338 0 57.0000pH 
K338 Lg338 Lflux338 1

Cg338 675 0 50.0000fF 
Lg338 675 676 57.0000pH
B338 675 676 10337 jj0 
Cgg338 676 0 50.0000fF
Vmeas338 676 677 0V

*Flux Biasing 
Idc339 0 50339 pwl(0 0uA 5ns 14.0680uA) 
Lflux339 50339 0 57.0000pH 
K339 Lg339 Lflux339 1

Cg339 677 0 50.0000fF 
Lg339 677 678 57.0000pH
B339 677 678 10338 jj0 
Cgg339 678 0 50.0000fF
Vmeas339 678 679 0V

*Flux Biasing 
Idc340 0 50340 pwl(0 0uA 5ns 14.0680uA) 
Lflux340 50340 0 57.0000pH 
K340 Lg340 Lflux340 1

Cg340 679 0 50.0000fF 
Lg340 679 680 57.0000pH
B340 679 680 10339 jj0 
Cgg340 680 0 50.0000fF
Vmeas340 680 681 0V

*Flux Biasing 
Idc341 0 50341 pwl(0 0uA 5ns 14.0680uA) 
Lflux341 50341 0 57.0000pH 
K341 Lg341 Lflux341 1

Cg341 681 0 50.0000fF 
Lg341 681 682 57.0000pH
B341 681 682 10340 jj0 
Cgg341 682 0 50.0000fF
Vmeas341 682 683 0V

*Flux Biasing 
Idc342 0 50342 pwl(0 0uA 5ns 14.0680uA) 
Lflux342 50342 0 57.0000pH 
K342 Lg342 Lflux342 1

Cg342 683 0 50.0000fF 
Lg342 683 684 57.0000pH
B342 683 684 10341 jj0 
Cgg342 684 0 50.0000fF
Vmeas342 684 685 0V

*Flux Biasing 
Idc343 0 50343 pwl(0 0uA 5ns 14.0680uA) 
Lflux343 50343 0 57.0000pH 
K343 Lg343 Lflux343 1

Cg343 685 0 50.0000fF 
Lg343 685 686 57.0000pH
B343 685 686 10342 jj0 
Cgg343 686 0 50.0000fF
Vmeas343 686 687 0V

*Flux Biasing 
Idc344 0 50344 pwl(0 0uA 5ns 14.0680uA) 
Lflux344 50344 0 57.0000pH 
K344 Lg344 Lflux344 1

Cg344 687 0 50.0000fF 
Lg344 687 688 57.0000pH
B344 687 688 10343 jj0 
Cgg344 688 0 50.0000fF
Vmeas344 688 689 0V

*Flux Biasing 
Idc345 0 50345 pwl(0 0uA 5ns 14.0680uA) 
Lflux345 50345 0 57.0000pH 
K345 Lg345 Lflux345 1

Cg345 689 0 50.0000fF 
Lg345 689 690 57.0000pH
B345 689 690 10344 jj0 
Cgg345 690 0 50.0000fF
Vmeas345 690 691 0V

*Flux Biasing 
Idc346 0 50346 pwl(0 0uA 5ns 14.0680uA) 
Lflux346 50346 0 57.0000pH 
K346 Lg346 Lflux346 1

Cg346 691 0 50.0000fF 
Lg346 691 692 57.0000pH
B346 691 692 10345 jj0 
Cgg346 692 0 50.0000fF
Vmeas346 692 693 0V

*Flux Biasing 
Idc347 0 50347 pwl(0 0uA 5ns 14.0680uA) 
Lflux347 50347 0 57.0000pH 
K347 Lg347 Lflux347 1

Cg347 693 0 50.0000fF 
Lg347 693 694 57.0000pH
B347 693 694 10346 jj0 
Cgg347 694 0 50.0000fF
Vmeas347 694 695 0V

*Flux Biasing 
Idc348 0 50348 pwl(0 0uA 5ns 14.0680uA) 
Lflux348 50348 0 57.0000pH 
K348 Lg348 Lflux348 1

Cg348 695 0 50.0000fF 
Lg348 695 696 57.0000pH
B348 695 696 10347 jj0 
Cgg348 696 0 50.0000fF
Vmeas348 696 697 0V

*Flux Biasing 
Idc349 0 50349 pwl(0 0uA 5ns 14.0680uA) 
Lflux349 50349 0 57.0000pH 
K349 Lg349 Lflux349 1

Cg349 697 0 50.0000fF 
Lg349 697 698 57.0000pH
B349 697 698 10348 jj0 
Cgg349 698 0 50.0000fF
Vmeas349 698 699 0V

*Flux Biasing 
Idc350 0 50350 pwl(0 0uA 5ns 14.0680uA) 
Lflux350 50350 0 57.0000pH 
K350 Lg350 Lflux350 1

Cg350 699 0 50.0000fF 
Lg350 699 700 57.0000pH
B350 699 700 10349 jj0 
Cgg350 700 0 50.0000fF
Vmeas350 700 701 0V

*Flux Biasing 
Idc351 0 50351 pwl(0 0uA 5ns 14.0680uA) 
Lflux351 50351 0 57.0000pH 
K351 Lg351 Lflux351 1

Cg351 701 0 50.0000fF 
Lg351 701 702 57.0000pH
B351 701 702 10350 jj0 
Cgg351 702 0 50.0000fF
Vmeas351 702 703 0V

*Flux Biasing 
Idc352 0 50352 pwl(0 0uA 5ns 14.0680uA) 
Lflux352 50352 0 57.0000pH 
K352 Lg352 Lflux352 1

Cg352 703 0 50.0000fF 
Lg352 703 704 57.0000pH
B352 703 704 10351 jj0 
Cgg352 704 0 50.0000fF
Vmeas352 704 705 0V

*Flux Biasing 
Idc353 0 50353 pwl(0 0uA 5ns 14.0680uA) 
Lflux353 50353 0 57.0000pH 
K353 Lg353 Lflux353 1

Cg353 705 0 50.0000fF 
Lg353 705 706 57.0000pH
B353 705 706 10352 jj0 
Cgg353 706 0 50.0000fF
Vmeas353 706 707 0V

*Flux Biasing 
Idc354 0 50354 pwl(0 0uA 5ns 14.0680uA) 
Lflux354 50354 0 57.0000pH 
K354 Lg354 Lflux354 1

Cg354 707 0 50.0000fF 
Lg354 707 708 57.0000pH
B354 707 708 10353 jj0 
Cgg354 708 0 50.0000fF
Vmeas354 708 709 0V

*Flux Biasing 
Idc355 0 50355 pwl(0 0uA 5ns 14.0680uA) 
Lflux355 50355 0 57.0000pH 
K355 Lg355 Lflux355 1

Cg355 709 0 50.0000fF 
Lg355 709 710 57.0000pH
B355 709 710 10354 jj0 
Cgg355 710 0 50.0000fF
Vmeas355 710 711 0V

*Flux Biasing 
Idc356 0 50356 pwl(0 0uA 5ns 14.0680uA) 
Lflux356 50356 0 57.0000pH 
K356 Lg356 Lflux356 1

Cg356 711 0 50.0000fF 
Lg356 711 712 57.0000pH
B356 711 712 10355 jj0 
Cgg356 712 0 50.0000fF
Vmeas356 712 713 0V

*Flux Biasing 
Idc357 0 50357 pwl(0 0uA 5ns 14.0680uA) 
Lflux357 50357 0 57.0000pH 
K357 Lg357 Lflux357 1

Cg357 713 0 50.0000fF 
Lg357 713 714 57.0000pH
B357 713 714 10356 jj0 
Cgg357 714 0 50.0000fF
Vmeas357 714 715 0V

*Flux Biasing 
Idc358 0 50358 pwl(0 0uA 5ns 14.0680uA) 
Lflux358 50358 0 57.0000pH 
K358 Lg358 Lflux358 1

Cg358 715 0 50.0000fF 
Lg358 715 716 57.0000pH
B358 715 716 10357 jj0 
Cgg358 716 0 50.0000fF
Vmeas358 716 717 0V

*Flux Biasing 
Idc359 0 50359 pwl(0 0uA 5ns 14.0680uA) 
Lflux359 50359 0 57.0000pH 
K359 Lg359 Lflux359 1

Cg359 717 0 50.0000fF 
Lg359 717 718 57.0000pH
B359 717 718 10358 jj0 
Cgg359 718 0 50.0000fF
Vmeas359 718 719 0V

*Flux Biasing 
Idc360 0 50360 pwl(0 0uA 5ns 14.0680uA) 
Lflux360 50360 0 57.0000pH 
K360 Lg360 Lflux360 1

Cg360 719 0 50.0000fF 
Lg360 719 720 57.0000pH
B360 719 720 10359 jj0 
Cgg360 720 0 50.0000fF
Vmeas360 720 721 0V

*Flux Biasing 
Idc361 0 50361 pwl(0 0uA 5ns 14.0680uA) 
Lflux361 50361 0 57.0000pH 
K361 Lg361 Lflux361 1

Cg361 721 0 50.0000fF 
Lg361 721 722 57.0000pH
B361 721 722 10360 jj0 
Cgg361 722 0 50.0000fF
Vmeas361 722 723 0V

*Flux Biasing 
Idc362 0 50362 pwl(0 0uA 5ns 14.0680uA) 
Lflux362 50362 0 57.0000pH 
K362 Lg362 Lflux362 1

Cg362 723 0 50.0000fF 
Lg362 723 724 57.0000pH
B362 723 724 10361 jj0 
Cgg362 724 0 50.0000fF
Vmeas362 724 725 0V

*Flux Biasing 
Idc363 0 50363 pwl(0 0uA 5ns 14.0680uA) 
Lflux363 50363 0 57.0000pH 
K363 Lg363 Lflux363 1

Cg363 725 0 50.0000fF 
Lg363 725 726 57.0000pH
B363 725 726 10362 jj0 
Cgg363 726 0 50.0000fF
Vmeas363 726 727 0V

*Flux Biasing 
Idc364 0 50364 pwl(0 0uA 5ns 14.0680uA) 
Lflux364 50364 0 57.0000pH 
K364 Lg364 Lflux364 1

Cg364 727 0 50.0000fF 
Lg364 727 728 57.0000pH
B364 727 728 10363 jj0 
Cgg364 728 0 50.0000fF
Vmeas364 728 729 0V

*Flux Biasing 
Idc365 0 50365 pwl(0 0uA 5ns 14.0680uA) 
Lflux365 50365 0 57.0000pH 
K365 Lg365 Lflux365 1

Cg365 729 0 50.0000fF 
Lg365 729 730 57.0000pH
B365 729 730 10364 jj0 
Cgg365 730 0 50.0000fF
Vmeas365 730 731 0V

*Flux Biasing 
Idc366 0 50366 pwl(0 0uA 5ns 14.0680uA) 
Lflux366 50366 0 57.0000pH 
K366 Lg366 Lflux366 1

Cg366 731 0 50.0000fF 
Lg366 731 732 57.0000pH
B366 731 732 10365 jj0 
Cgg366 732 0 50.0000fF
Vmeas366 732 733 0V

*Flux Biasing 
Idc367 0 50367 pwl(0 0uA 5ns 14.0680uA) 
Lflux367 50367 0 57.0000pH 
K367 Lg367 Lflux367 1

Cg367 733 0 50.0000fF 
Lg367 733 734 57.0000pH
B367 733 734 10366 jj0 
Cgg367 734 0 50.0000fF
Vmeas367 734 735 0V

*Flux Biasing 
Idc368 0 50368 pwl(0 0uA 5ns 14.0680uA) 
Lflux368 50368 0 57.0000pH 
K368 Lg368 Lflux368 1

Cg368 735 0 50.0000fF 
Lg368 735 736 57.0000pH
B368 735 736 10367 jj0 
Cgg368 736 0 50.0000fF
Vmeas368 736 737 0V

*Flux Biasing 
Idc369 0 50369 pwl(0 0uA 5ns 14.0680uA) 
Lflux369 50369 0 57.0000pH 
K369 Lg369 Lflux369 1

Cg369 737 0 50.0000fF 
Lg369 737 738 57.0000pH
B369 737 738 10368 jj0 
Cgg369 738 0 50.0000fF
Vmeas369 738 739 0V

*Flux Biasing 
Idc370 0 50370 pwl(0 0uA 5ns 14.0680uA) 
Lflux370 50370 0 57.0000pH 
K370 Lg370 Lflux370 1

Cg370 739 0 50.0000fF 
Lg370 739 740 57.0000pH
B370 739 740 10369 jj0 
Cgg370 740 0 50.0000fF
Vmeas370 740 741 0V

*Flux Biasing 
Idc371 0 50371 pwl(0 0uA 5ns 14.0680uA) 
Lflux371 50371 0 57.0000pH 
K371 Lg371 Lflux371 1

Cg371 741 0 50.0000fF 
Lg371 741 742 57.0000pH
B371 741 742 10370 jj0 
Cgg371 742 0 50.0000fF
Vmeas371 742 743 0V

*Flux Biasing 
Idc372 0 50372 pwl(0 0uA 5ns 14.0680uA) 
Lflux372 50372 0 57.0000pH 
K372 Lg372 Lflux372 1

Cg372 743 0 50.0000fF 
Lg372 743 744 57.0000pH
B372 743 744 10371 jj0 
Cgg372 744 0 50.0000fF
Vmeas372 744 745 0V

*Flux Biasing 
Idc373 0 50373 pwl(0 0uA 5ns 14.0680uA) 
Lflux373 50373 0 57.0000pH 
K373 Lg373 Lflux373 1

Cg373 745 0 50.0000fF 
Lg373 745 746 57.0000pH
B373 745 746 10372 jj0 
Cgg373 746 0 50.0000fF
Vmeas373 746 747 0V

*Flux Biasing 
Idc374 0 50374 pwl(0 0uA 5ns 14.0680uA) 
Lflux374 50374 0 57.0000pH 
K374 Lg374 Lflux374 1

Cg374 747 0 50.0000fF 
Lg374 747 748 57.0000pH
B374 747 748 10373 jj0 
Cgg374 748 0 50.0000fF
Vmeas374 748 749 0V

*Flux Biasing 
Idc375 0 50375 pwl(0 0uA 5ns 14.0680uA) 
Lflux375 50375 0 57.0000pH 
K375 Lg375 Lflux375 1

Cg375 749 0 50.0000fF 
Lg375 749 750 57.0000pH
B375 749 750 10374 jj0 
Cgg375 750 0 50.0000fF
Vmeas375 750 751 0V

*Flux Biasing 
Idc376 0 50376 pwl(0 0uA 5ns 14.0680uA) 
Lflux376 50376 0 57.0000pH 
K376 Lg376 Lflux376 1

Cg376 751 0 50.0000fF 
Lg376 751 752 57.0000pH
B376 751 752 10375 jj0 
Cgg376 752 0 50.0000fF
Vmeas376 752 753 0V

*Flux Biasing 
Idc377 0 50377 pwl(0 0uA 5ns 14.0680uA) 
Lflux377 50377 0 57.0000pH 
K377 Lg377 Lflux377 1

Cg377 753 0 50.0000fF 
Lg377 753 754 57.0000pH
B377 753 754 10376 jj0 
Cgg377 754 0 50.0000fF
Vmeas377 754 755 0V

*Flux Biasing 
Idc378 0 50378 pwl(0 0uA 5ns 14.0680uA) 
Lflux378 50378 0 57.0000pH 
K378 Lg378 Lflux378 1

Cg378 755 0 50.0000fF 
Lg378 755 756 57.0000pH
B378 755 756 10377 jj0 
Cgg378 756 0 50.0000fF
Vmeas378 756 757 0V

*Flux Biasing 
Idc379 0 50379 pwl(0 0uA 5ns 14.0680uA) 
Lflux379 50379 0 57.0000pH 
K379 Lg379 Lflux379 1

Cg379 757 0 50.0000fF 
Lg379 757 758 57.0000pH
B379 757 758 10378 jj0 
Cgg379 758 0 50.0000fF
Vmeas379 758 759 0V

*Flux Biasing 
Idc380 0 50380 pwl(0 0uA 5ns 14.0680uA) 
Lflux380 50380 0 57.0000pH 
K380 Lg380 Lflux380 1

Cg380 759 0 50.0000fF 
Lg380 759 760 57.0000pH
B380 759 760 10379 jj0 
Cgg380 760 0 50.0000fF
Vmeas380 760 761 0V

*Flux Biasing 
Idc381 0 50381 pwl(0 0uA 5ns 14.0680uA) 
Lflux381 50381 0 57.0000pH 
K381 Lg381 Lflux381 1

Cg381 761 0 50.0000fF 
Lg381 761 762 57.0000pH
B381 761 762 10380 jj0 
Cgg381 762 0 50.0000fF
Vmeas381 762 763 0V

*Flux Biasing 
Idc382 0 50382 pwl(0 0uA 5ns 14.0680uA) 
Lflux382 50382 0 57.0000pH 
K382 Lg382 Lflux382 1

Cg382 763 0 50.0000fF 
Lg382 763 764 57.0000pH
B382 763 764 10381 jj0 
Cgg382 764 0 50.0000fF
Vmeas382 764 765 0V

*Flux Biasing 
Idc383 0 50383 pwl(0 0uA 5ns 14.0680uA) 
Lflux383 50383 0 57.0000pH 
K383 Lg383 Lflux383 1

Cg383 765 0 50.0000fF 
Lg383 765 766 57.0000pH
B383 765 766 10382 jj0 
Cgg383 766 0 50.0000fF
Vmeas383 766 767 0V

*Flux Biasing 
Idc384 0 50384 pwl(0 0uA 5ns 14.0680uA) 
Lflux384 50384 0 57.0000pH 
K384 Lg384 Lflux384 1

Cg384 767 0 50.0000fF 
Lg384 767 768 57.0000pH
B384 767 768 10383 jj0 
Cgg384 768 0 50.0000fF
Vmeas384 768 769 0V

*Flux Biasing 
Idc385 0 50385 pwl(0 0uA 5ns 14.0680uA) 
Lflux385 50385 0 57.0000pH 
K385 Lg385 Lflux385 1

Cg385 769 0 50.0000fF 
Lg385 769 770 57.0000pH
B385 769 770 10384 jj0 
Cgg385 770 0 50.0000fF
Vmeas385 770 771 0V

*Flux Biasing 
Idc386 0 50386 pwl(0 0uA 5ns 14.0680uA) 
Lflux386 50386 0 57.0000pH 
K386 Lg386 Lflux386 1

Cg386 771 0 50.0000fF 
Lg386 771 772 57.0000pH
B386 771 772 10385 jj0 
Cgg386 772 0 50.0000fF
Vmeas386 772 773 0V

*Flux Biasing 
Idc387 0 50387 pwl(0 0uA 5ns 14.0680uA) 
Lflux387 50387 0 57.0000pH 
K387 Lg387 Lflux387 1

Cg387 773 0 50.0000fF 
Lg387 773 774 57.0000pH
B387 773 774 10386 jj0 
Cgg387 774 0 50.0000fF
Vmeas387 774 775 0V

*Flux Biasing 
Idc388 0 50388 pwl(0 0uA 5ns 14.0680uA) 
Lflux388 50388 0 57.0000pH 
K388 Lg388 Lflux388 1

Cg388 775 0 50.0000fF 
Lg388 775 776 57.0000pH
B388 775 776 10387 jj0 
Cgg388 776 0 50.0000fF
Vmeas388 776 777 0V

*Flux Biasing 
Idc389 0 50389 pwl(0 0uA 5ns 14.0680uA) 
Lflux389 50389 0 57.0000pH 
K389 Lg389 Lflux389 1

Cg389 777 0 50.0000fF 
Lg389 777 778 57.0000pH
B389 777 778 10388 jj0 
Cgg389 778 0 50.0000fF
Vmeas389 778 779 0V

*Flux Biasing 
Idc390 0 50390 pwl(0 0uA 5ns 14.0680uA) 
Lflux390 50390 0 57.0000pH 
K390 Lg390 Lflux390 1

Cg390 779 0 50.0000fF 
Lg390 779 780 57.0000pH
B390 779 780 10389 jj0 
Cgg390 780 0 50.0000fF
Vmeas390 780 781 0V

*Flux Biasing 
Idc391 0 50391 pwl(0 0uA 5ns 14.0680uA) 
Lflux391 50391 0 57.0000pH 
K391 Lg391 Lflux391 1

Cg391 781 0 50.0000fF 
Lg391 781 782 57.0000pH
B391 781 782 10390 jj0 
Cgg391 782 0 50.0000fF
Vmeas391 782 783 0V

*Flux Biasing 
Idc392 0 50392 pwl(0 0uA 5ns 14.0680uA) 
Lflux392 50392 0 57.0000pH 
K392 Lg392 Lflux392 1

Cg392 783 0 50.0000fF 
Lg392 783 784 57.0000pH
B392 783 784 10391 jj0 
Cgg392 784 0 50.0000fF
Vmeas392 784 785 0V

*Flux Biasing 
Idc393 0 50393 pwl(0 0uA 5ns 14.0680uA) 
Lflux393 50393 0 57.0000pH 
K393 Lg393 Lflux393 1

Cg393 785 0 50.0000fF 
Lg393 785 786 57.0000pH
B393 785 786 10392 jj0 
Cgg393 786 0 50.0000fF
Vmeas393 786 787 0V

*Flux Biasing 
Idc394 0 50394 pwl(0 0uA 5ns 14.0680uA) 
Lflux394 50394 0 57.0000pH 
K394 Lg394 Lflux394 1

Cg394 787 0 50.0000fF 
Lg394 787 788 57.0000pH
B394 787 788 10393 jj0 
Cgg394 788 0 50.0000fF
Vmeas394 788 789 0V

*Flux Biasing 
Idc395 0 50395 pwl(0 0uA 5ns 14.0680uA) 
Lflux395 50395 0 57.0000pH 
K395 Lg395 Lflux395 1

Cg395 789 0 50.0000fF 
Lg395 789 790 57.0000pH
B395 789 790 10394 jj0 
Cgg395 790 0 50.0000fF
Vmeas395 790 791 0V

*Flux Biasing 
Idc396 0 50396 pwl(0 0uA 5ns 14.0680uA) 
Lflux396 50396 0 57.0000pH 
K396 Lg396 Lflux396 1

Cg396 791 0 50.0000fF 
Lg396 791 792 57.0000pH
B396 791 792 10395 jj0 
Cgg396 792 0 50.0000fF
Vmeas396 792 793 0V

*Flux Biasing 
Idc397 0 50397 pwl(0 0uA 5ns 14.0680uA) 
Lflux397 50397 0 57.0000pH 
K397 Lg397 Lflux397 1

Cg397 793 0 50.0000fF 
Lg397 793 794 57.0000pH
B397 793 794 10396 jj0 
Cgg397 794 0 50.0000fF
Vmeas397 794 795 0V

*Flux Biasing 
Idc398 0 50398 pwl(0 0uA 5ns 14.0680uA) 
Lflux398 50398 0 57.0000pH 
K398 Lg398 Lflux398 1

Cg398 795 0 50.0000fF 
Lg398 795 796 57.0000pH
B398 795 796 10397 jj0 
Cgg398 796 0 50.0000fF
Vmeas398 796 797 0V

*Flux Biasing 
Idc399 0 50399 pwl(0 0uA 5ns 14.0680uA) 
Lflux399 50399 0 57.0000pH 
K399 Lg399 Lflux399 1

Cg399 797 0 50.0000fF 
Lg399 797 798 57.0000pH
B399 797 798 10398 jj0 
Cgg399 798 0 50.0000fF
Vmeas399 798 799 0V

*Flux Biasing 
Idc400 0 50400 pwl(0 0uA 5ns 14.0680uA) 
Lflux400 50400 0 57.0000pH 
K400 Lg400 Lflux400 1

Cg400 799 0 50.0000fF 
Lg400 799 800 57.0000pH
B400 799 800 10399 jj0 
Cgg400 800 0 50.0000fF
Vmeas400 800 801 0V

*Flux Biasing 
Idc401 0 50401 pwl(0 0uA 5ns 14.0680uA) 
Lflux401 50401 0 57.0000pH 
K401 Lg401 Lflux401 1

Cg401 801 0 50.0000fF 
Lg401 801 802 57.0000pH
B401 801 802 10400 jj0 
Cgg401 802 0 50.0000fF
Vmeas401 802 803 0V

*Flux Biasing 
Idc402 0 50402 pwl(0 0uA 5ns 14.0680uA) 
Lflux402 50402 0 57.0000pH 
K402 Lg402 Lflux402 1

Cg402 803 0 50.0000fF 
Lg402 803 804 57.0000pH
B402 803 804 10401 jj0 
Cgg402 804 0 50.0000fF
Vmeas402 804 805 0V

*Flux Biasing 
Idc403 0 50403 pwl(0 0uA 5ns 14.0680uA) 
Lflux403 50403 0 57.0000pH 
K403 Lg403 Lflux403 1

Cg403 805 0 50.0000fF 
Lg403 805 806 57.0000pH
B403 805 806 10402 jj0 
Cgg403 806 0 50.0000fF
Vmeas403 806 807 0V

*Flux Biasing 
Idc404 0 50404 pwl(0 0uA 5ns 14.0680uA) 
Lflux404 50404 0 57.0000pH 
K404 Lg404 Lflux404 1

Cg404 807 0 50.0000fF 
Lg404 807 808 57.0000pH
B404 807 808 10403 jj0 
Cgg404 808 0 50.0000fF
Vmeas404 808 809 0V

*Flux Biasing 
Idc405 0 50405 pwl(0 0uA 5ns 14.0680uA) 
Lflux405 50405 0 57.0000pH 
K405 Lg405 Lflux405 1

Cg405 809 0 50.0000fF 
Lg405 809 810 57.0000pH
B405 809 810 10404 jj0 
Cgg405 810 0 50.0000fF
Vmeas405 810 811 0V

*Flux Biasing 
Idc406 0 50406 pwl(0 0uA 5ns 14.0680uA) 
Lflux406 50406 0 57.0000pH 
K406 Lg406 Lflux406 1

Cg406 811 0 50.0000fF 
Lg406 811 812 57.0000pH
B406 811 812 10405 jj0 
Cgg406 812 0 50.0000fF
Vmeas406 812 813 0V

*Flux Biasing 
Idc407 0 50407 pwl(0 0uA 5ns 14.0680uA) 
Lflux407 50407 0 57.0000pH 
K407 Lg407 Lflux407 1

Cg407 813 0 50.0000fF 
Lg407 813 814 57.0000pH
B407 813 814 10406 jj0 
Cgg407 814 0 50.0000fF
Vmeas407 814 815 0V

*Flux Biasing 
Idc408 0 50408 pwl(0 0uA 5ns 14.0680uA) 
Lflux408 50408 0 57.0000pH 
K408 Lg408 Lflux408 1

Cg408 815 0 50.0000fF 
Lg408 815 816 57.0000pH
B408 815 816 10407 jj0 
Cgg408 816 0 50.0000fF
Vmeas408 816 817 0V

*Flux Biasing 
Idc409 0 50409 pwl(0 0uA 5ns 14.0680uA) 
Lflux409 50409 0 57.0000pH 
K409 Lg409 Lflux409 1

Cg409 817 0 50.0000fF 
Lg409 817 818 57.0000pH
B409 817 818 10408 jj0 
Cgg409 818 0 50.0000fF
Vmeas409 818 819 0V

*Flux Biasing 
Idc410 0 50410 pwl(0 0uA 5ns 14.0680uA) 
Lflux410 50410 0 57.0000pH 
K410 Lg410 Lflux410 1

Cg410 819 0 50.0000fF 
Lg410 819 820 57.0000pH
B410 819 820 10409 jj0 
Cgg410 820 0 50.0000fF
Vmeas410 820 821 0V

*Flux Biasing 
Idc411 0 50411 pwl(0 0uA 5ns 14.0680uA) 
Lflux411 50411 0 57.0000pH 
K411 Lg411 Lflux411 1

Cg411 821 0 50.0000fF 
Lg411 821 822 57.0000pH
B411 821 822 10410 jj0 
Cgg411 822 0 50.0000fF
Vmeas411 822 823 0V

*Flux Biasing 
Idc412 0 50412 pwl(0 0uA 5ns 14.0680uA) 
Lflux412 50412 0 57.0000pH 
K412 Lg412 Lflux412 1

Cg412 823 0 50.0000fF 
Lg412 823 824 57.0000pH
B412 823 824 10411 jj0 
Cgg412 824 0 50.0000fF
Vmeas412 824 825 0V

*Flux Biasing 
Idc413 0 50413 pwl(0 0uA 5ns 14.0680uA) 
Lflux413 50413 0 57.0000pH 
K413 Lg413 Lflux413 1

Cg413 825 0 50.0000fF 
Lg413 825 826 57.0000pH
B413 825 826 10412 jj0 
Cgg413 826 0 50.0000fF
Vmeas413 826 827 0V

*Flux Biasing 
Idc414 0 50414 pwl(0 0uA 5ns 14.0680uA) 
Lflux414 50414 0 57.0000pH 
K414 Lg414 Lflux414 1

Cg414 827 0 50.0000fF 
Lg414 827 828 57.0000pH
B414 827 828 10413 jj0 
Cgg414 828 0 50.0000fF
Vmeas414 828 829 0V

*Flux Biasing 
Idc415 0 50415 pwl(0 0uA 5ns 14.0680uA) 
Lflux415 50415 0 57.0000pH 
K415 Lg415 Lflux415 1

Cg415 829 0 50.0000fF 
Lg415 829 830 57.0000pH
B415 829 830 10414 jj0 
Cgg415 830 0 50.0000fF
Vmeas415 830 831 0V

*Flux Biasing 
Idc416 0 50416 pwl(0 0uA 5ns 14.0680uA) 
Lflux416 50416 0 57.0000pH 
K416 Lg416 Lflux416 1

Cg416 831 0 50.0000fF 
Lg416 831 832 57.0000pH
B416 831 832 10415 jj0 
Cgg416 832 0 50.0000fF
Vmeas416 832 833 0V

*Flux Biasing 
Idc417 0 50417 pwl(0 0uA 5ns 14.0680uA) 
Lflux417 50417 0 57.0000pH 
K417 Lg417 Lflux417 1

Cg417 833 0 50.0000fF 
Lg417 833 834 57.0000pH
B417 833 834 10416 jj0 
Cgg417 834 0 50.0000fF
Vmeas417 834 835 0V

*Flux Biasing 
Idc418 0 50418 pwl(0 0uA 5ns 14.0680uA) 
Lflux418 50418 0 57.0000pH 
K418 Lg418 Lflux418 1

Cg418 835 0 50.0000fF 
Lg418 835 836 57.0000pH
B418 835 836 10417 jj0 
Cgg418 836 0 50.0000fF
Vmeas418 836 837 0V

*Flux Biasing 
Idc419 0 50419 pwl(0 0uA 5ns 14.0680uA) 
Lflux419 50419 0 57.0000pH 
K419 Lg419 Lflux419 1

Cg419 837 0 50.0000fF 
Lg419 837 838 57.0000pH
B419 837 838 10418 jj0 
Cgg419 838 0 50.0000fF
Vmeas419 838 839 0V

*Flux Biasing 
Idc420 0 50420 pwl(0 0uA 5ns 14.0680uA) 
Lflux420 50420 0 57.0000pH 
K420 Lg420 Lflux420 1

Cg420 839 0 50.0000fF 
Lg420 839 840 57.0000pH
B420 839 840 10419 jj0 
Cgg420 840 0 50.0000fF
Vmeas420 840 841 0V

*Flux Biasing 
Idc421 0 50421 pwl(0 0uA 5ns 14.0680uA) 
Lflux421 50421 0 57.0000pH 
K421 Lg421 Lflux421 1

Cg421 841 0 50.0000fF 
Lg421 841 842 57.0000pH
B421 841 842 10420 jj0 
Cgg421 842 0 50.0000fF
Vmeas421 842 843 0V

*Flux Biasing 
Idc422 0 50422 pwl(0 0uA 5ns 14.0680uA) 
Lflux422 50422 0 57.0000pH 
K422 Lg422 Lflux422 1

Cg422 843 0 50.0000fF 
Lg422 843 844 57.0000pH
B422 843 844 10421 jj0 
Cgg422 844 0 50.0000fF
Vmeas422 844 845 0V

*Flux Biasing 
Idc423 0 50423 pwl(0 0uA 5ns 14.0680uA) 
Lflux423 50423 0 57.0000pH 
K423 Lg423 Lflux423 1

Cg423 845 0 50.0000fF 
Lg423 845 846 57.0000pH
B423 845 846 10422 jj0 
Cgg423 846 0 50.0000fF
Vmeas423 846 847 0V

*Flux Biasing 
Idc424 0 50424 pwl(0 0uA 5ns 14.0680uA) 
Lflux424 50424 0 57.0000pH 
K424 Lg424 Lflux424 1

Cg424 847 0 50.0000fF 
Lg424 847 848 57.0000pH
B424 847 848 10423 jj0 
Cgg424 848 0 50.0000fF
Vmeas424 848 849 0V

*Flux Biasing 
Idc425 0 50425 pwl(0 0uA 5ns 14.0680uA) 
Lflux425 50425 0 57.0000pH 
K425 Lg425 Lflux425 1

Cg425 849 0 50.0000fF 
Lg425 849 850 57.0000pH
B425 849 850 10424 jj0 
Cgg425 850 0 50.0000fF
Vmeas425 850 851 0V

*Flux Biasing 
Idc426 0 50426 pwl(0 0uA 5ns 14.0680uA) 
Lflux426 50426 0 57.0000pH 
K426 Lg426 Lflux426 1

Cg426 851 0 50.0000fF 
Lg426 851 852 57.0000pH
B426 851 852 10425 jj0 
Cgg426 852 0 50.0000fF
Vmeas426 852 853 0V

*Flux Biasing 
Idc427 0 50427 pwl(0 0uA 5ns 14.0680uA) 
Lflux427 50427 0 57.0000pH 
K427 Lg427 Lflux427 1

Cg427 853 0 50.0000fF 
Lg427 853 854 57.0000pH
B427 853 854 10426 jj0 
Cgg427 854 0 50.0000fF
Vmeas427 854 855 0V

*Flux Biasing 
Idc428 0 50428 pwl(0 0uA 5ns 14.0680uA) 
Lflux428 50428 0 57.0000pH 
K428 Lg428 Lflux428 1

Cg428 855 0 50.0000fF 
Lg428 855 856 57.0000pH
B428 855 856 10427 jj0 
Cgg428 856 0 50.0000fF
Vmeas428 856 857 0V

*Flux Biasing 
Idc429 0 50429 pwl(0 0uA 5ns 14.0680uA) 
Lflux429 50429 0 57.0000pH 
K429 Lg429 Lflux429 1

Cg429 857 0 50.0000fF 
Lg429 857 858 57.0000pH
B429 857 858 10428 jj0 
Cgg429 858 0 50.0000fF
Vmeas429 858 859 0V

*Flux Biasing 
Idc430 0 50430 pwl(0 0uA 5ns 14.0680uA) 
Lflux430 50430 0 57.0000pH 
K430 Lg430 Lflux430 1

Cg430 859 0 50.0000fF 
Lg430 859 860 57.0000pH
B430 859 860 10429 jj0 
Cgg430 860 0 50.0000fF
Vmeas430 860 861 0V

*Flux Biasing 
Idc431 0 50431 pwl(0 0uA 5ns 14.0680uA) 
Lflux431 50431 0 57.0000pH 
K431 Lg431 Lflux431 1

Cg431 861 0 50.0000fF 
Lg431 861 862 57.0000pH
B431 861 862 10430 jj0 
Cgg431 862 0 50.0000fF
Vmeas431 862 863 0V

*Flux Biasing 
Idc432 0 50432 pwl(0 0uA 5ns 14.0680uA) 
Lflux432 50432 0 57.0000pH 
K432 Lg432 Lflux432 1

Cg432 863 0 50.0000fF 
Lg432 863 864 57.0000pH
B432 863 864 10431 jj0 
Cgg432 864 0 50.0000fF
Vmeas432 864 865 0V

*Flux Biasing 
Idc433 0 50433 pwl(0 0uA 5ns 14.0680uA) 
Lflux433 50433 0 57.0000pH 
K433 Lg433 Lflux433 1

Cg433 865 0 50.0000fF 
Lg433 865 866 57.0000pH
B433 865 866 10432 jj0 
Cgg433 866 0 50.0000fF
Vmeas433 866 867 0V

*Flux Biasing 
Idc434 0 50434 pwl(0 0uA 5ns 14.0680uA) 
Lflux434 50434 0 57.0000pH 
K434 Lg434 Lflux434 1

Cg434 867 0 50.0000fF 
Lg434 867 868 57.0000pH
B434 867 868 10433 jj0 
Cgg434 868 0 50.0000fF
Vmeas434 868 869 0V

*Flux Biasing 
Idc435 0 50435 pwl(0 0uA 5ns 14.0680uA) 
Lflux435 50435 0 57.0000pH 
K435 Lg435 Lflux435 1

Cg435 869 0 50.0000fF 
Lg435 869 870 57.0000pH
B435 869 870 10434 jj0 
Cgg435 870 0 50.0000fF
Vmeas435 870 871 0V

*Flux Biasing 
Idc436 0 50436 pwl(0 0uA 5ns 14.0680uA) 
Lflux436 50436 0 57.0000pH 
K436 Lg436 Lflux436 1

Cg436 871 0 50.0000fF 
Lg436 871 872 57.0000pH
B436 871 872 10435 jj0 
Cgg436 872 0 50.0000fF
Vmeas436 872 873 0V

*Flux Biasing 
Idc437 0 50437 pwl(0 0uA 5ns 14.0680uA) 
Lflux437 50437 0 57.0000pH 
K437 Lg437 Lflux437 1

Cg437 873 0 50.0000fF 
Lg437 873 874 57.0000pH
B437 873 874 10436 jj0 
Cgg437 874 0 50.0000fF
Vmeas437 874 875 0V

*Flux Biasing 
Idc438 0 50438 pwl(0 0uA 5ns 14.0680uA) 
Lflux438 50438 0 57.0000pH 
K438 Lg438 Lflux438 1

Cg438 875 0 50.0000fF 
Lg438 875 876 57.0000pH
B438 875 876 10437 jj0 
Cgg438 876 0 50.0000fF
Vmeas438 876 877 0V

*Flux Biasing 
Idc439 0 50439 pwl(0 0uA 5ns 14.0680uA) 
Lflux439 50439 0 57.0000pH 
K439 Lg439 Lflux439 1

Cg439 877 0 50.0000fF 
Lg439 877 878 57.0000pH
B439 877 878 10438 jj0 
Cgg439 878 0 50.0000fF
Vmeas439 878 879 0V

*Flux Biasing 
Idc440 0 50440 pwl(0 0uA 5ns 14.0680uA) 
Lflux440 50440 0 57.0000pH 
K440 Lg440 Lflux440 1

Cg440 879 0 50.0000fF 
Lg440 879 880 57.0000pH
B440 879 880 10439 jj0 
Cgg440 880 0 50.0000fF
Vmeas440 880 881 0V

*Flux Biasing 
Idc441 0 50441 pwl(0 0uA 5ns 14.0680uA) 
Lflux441 50441 0 57.0000pH 
K441 Lg441 Lflux441 1

Cg441 881 0 50.0000fF 
Lg441 881 882 57.0000pH
B441 881 882 10440 jj0 
Cgg441 882 0 50.0000fF
Vmeas441 882 883 0V

*Flux Biasing 
Idc442 0 50442 pwl(0 0uA 5ns 14.0680uA) 
Lflux442 50442 0 57.0000pH 
K442 Lg442 Lflux442 1

Cg442 883 0 50.0000fF 
Lg442 883 884 57.0000pH
B442 883 884 10441 jj0 
Cgg442 884 0 50.0000fF
Vmeas442 884 885 0V

*Flux Biasing 
Idc443 0 50443 pwl(0 0uA 5ns 14.0680uA) 
Lflux443 50443 0 57.0000pH 
K443 Lg443 Lflux443 1

Cg443 885 0 50.0000fF 
Lg443 885 886 57.0000pH
B443 885 886 10442 jj0 
Cgg443 886 0 50.0000fF
Vmeas443 886 887 0V

*Flux Biasing 
Idc444 0 50444 pwl(0 0uA 5ns 14.0680uA) 
Lflux444 50444 0 57.0000pH 
K444 Lg444 Lflux444 1

Cg444 887 0 50.0000fF 
Lg444 887 888 57.0000pH
B444 887 888 10443 jj0 
Cgg444 888 0 50.0000fF
Vmeas444 888 889 0V

*Flux Biasing 
Idc445 0 50445 pwl(0 0uA 5ns 14.0680uA) 
Lflux445 50445 0 57.0000pH 
K445 Lg445 Lflux445 1

Cg445 889 0 50.0000fF 
Lg445 889 890 57.0000pH
B445 889 890 10444 jj0 
Cgg445 890 0 50.0000fF
Vmeas445 890 891 0V

*Flux Biasing 
Idc446 0 50446 pwl(0 0uA 5ns 14.0680uA) 
Lflux446 50446 0 57.0000pH 
K446 Lg446 Lflux446 1

Cg446 891 0 50.0000fF 
Lg446 891 892 57.0000pH
B446 891 892 10445 jj0 
Cgg446 892 0 50.0000fF
Vmeas446 892 893 0V

*Flux Biasing 
Idc447 0 50447 pwl(0 0uA 5ns 14.0680uA) 
Lflux447 50447 0 57.0000pH 
K447 Lg447 Lflux447 1

Cg447 893 0 50.0000fF 
Lg447 893 894 57.0000pH
B447 893 894 10446 jj0 
Cgg447 894 0 50.0000fF
Vmeas447 894 895 0V

*Flux Biasing 
Idc448 0 50448 pwl(0 0uA 5ns 14.0680uA) 
Lflux448 50448 0 57.0000pH 
K448 Lg448 Lflux448 1

Cg448 895 0 50.0000fF 
Lg448 895 896 57.0000pH
B448 895 896 10447 jj0 
Cgg448 896 0 50.0000fF
Vmeas448 896 897 0V

*Flux Biasing 
Idc449 0 50449 pwl(0 0uA 5ns 14.0680uA) 
Lflux449 50449 0 57.0000pH 
K449 Lg449 Lflux449 1

Cg449 897 0 50.0000fF 
Lg449 897 898 57.0000pH
B449 897 898 10448 jj0 
Cgg449 898 0 50.0000fF
Vmeas449 898 899 0V

*Flux Biasing 
Idc450 0 50450 pwl(0 0uA 5ns 14.0680uA) 
Lflux450 50450 0 57.0000pH 
K450 Lg450 Lflux450 1

Cg450 899 0 50.0000fF 
Lg450 899 900 57.0000pH
B450 899 900 10449 jj0 
Cgg450 900 0 50.0000fF
Vmeas450 900 901 0V

*Flux Biasing 
Idc451 0 50451 pwl(0 0uA 5ns 14.0680uA) 
Lflux451 50451 0 57.0000pH 
K451 Lg451 Lflux451 1

Cg451 901 0 50.0000fF 
Lg451 901 902 57.0000pH
B451 901 902 10450 jj0 
Cgg451 902 0 50.0000fF
Vmeas451 902 903 0V

*Flux Biasing 
Idc452 0 50452 pwl(0 0uA 5ns 14.0680uA) 
Lflux452 50452 0 57.0000pH 
K452 Lg452 Lflux452 1

Cg452 903 0 50.0000fF 
Lg452 903 904 57.0000pH
B452 903 904 10451 jj0 
Cgg452 904 0 50.0000fF
Vmeas452 904 905 0V

*Flux Biasing 
Idc453 0 50453 pwl(0 0uA 5ns 14.0680uA) 
Lflux453 50453 0 57.0000pH 
K453 Lg453 Lflux453 1

Cg453 905 0 50.0000fF 
Lg453 905 906 57.0000pH
B453 905 906 10452 jj0 
Cgg453 906 0 50.0000fF
Vmeas453 906 907 0V

*Flux Biasing 
Idc454 0 50454 pwl(0 0uA 5ns 14.0680uA) 
Lflux454 50454 0 57.0000pH 
K454 Lg454 Lflux454 1

Cg454 907 0 50.0000fF 
Lg454 907 908 57.0000pH
B454 907 908 10453 jj0 
Cgg454 908 0 50.0000fF
Vmeas454 908 909 0V

*Flux Biasing 
Idc455 0 50455 pwl(0 0uA 5ns 14.0680uA) 
Lflux455 50455 0 57.0000pH 
K455 Lg455 Lflux455 1

Cg455 909 0 50.0000fF 
Lg455 909 910 57.0000pH
B455 909 910 10454 jj0 
Cgg455 910 0 50.0000fF
Vmeas455 910 911 0V

*Flux Biasing 
Idc456 0 50456 pwl(0 0uA 5ns 14.0680uA) 
Lflux456 50456 0 57.0000pH 
K456 Lg456 Lflux456 1

Cg456 911 0 50.0000fF 
Lg456 911 912 57.0000pH
B456 911 912 10455 jj0 
Cgg456 912 0 50.0000fF
Vmeas456 912 913 0V

*Flux Biasing 
Idc457 0 50457 pwl(0 0uA 5ns 14.0680uA) 
Lflux457 50457 0 57.0000pH 
K457 Lg457 Lflux457 1

Cg457 913 0 50.0000fF 
Lg457 913 914 57.0000pH
B457 913 914 10456 jj0 
Cgg457 914 0 50.0000fF
Vmeas457 914 915 0V

*Flux Biasing 
Idc458 0 50458 pwl(0 0uA 5ns 14.0680uA) 
Lflux458 50458 0 57.0000pH 
K458 Lg458 Lflux458 1

Cg458 915 0 50.0000fF 
Lg458 915 916 57.0000pH
B458 915 916 10457 jj0 
Cgg458 916 0 50.0000fF
Vmeas458 916 917 0V

*Flux Biasing 
Idc459 0 50459 pwl(0 0uA 5ns 14.0680uA) 
Lflux459 50459 0 57.0000pH 
K459 Lg459 Lflux459 1

Cg459 917 0 50.0000fF 
Lg459 917 918 57.0000pH
B459 917 918 10458 jj0 
Cgg459 918 0 50.0000fF
Vmeas459 918 919 0V

*Flux Biasing 
Idc460 0 50460 pwl(0 0uA 5ns 14.0680uA) 
Lflux460 50460 0 57.0000pH 
K460 Lg460 Lflux460 1

Cg460 919 0 50.0000fF 
Lg460 919 920 57.0000pH
B460 919 920 10459 jj0 
Cgg460 920 0 50.0000fF
Vmeas460 920 921 0V

*Flux Biasing 
Idc461 0 50461 pwl(0 0uA 5ns 14.0680uA) 
Lflux461 50461 0 57.0000pH 
K461 Lg461 Lflux461 1

Cg461 921 0 50.0000fF 
Lg461 921 922 57.0000pH
B461 921 922 10460 jj0 
Cgg461 922 0 50.0000fF
Vmeas461 922 923 0V

*Flux Biasing 
Idc462 0 50462 pwl(0 0uA 5ns 14.0680uA) 
Lflux462 50462 0 57.0000pH 
K462 Lg462 Lflux462 1

Cg462 923 0 50.0000fF 
Lg462 923 924 57.0000pH
B462 923 924 10461 jj0 
Cgg462 924 0 50.0000fF
Vmeas462 924 925 0V

*Flux Biasing 
Idc463 0 50463 pwl(0 0uA 5ns 14.0680uA) 
Lflux463 50463 0 57.0000pH 
K463 Lg463 Lflux463 1

Cg463 925 0 50.0000fF 
Lg463 925 926 57.0000pH
B463 925 926 10462 jj0 
Cgg463 926 0 50.0000fF
Vmeas463 926 927 0V

*Flux Biasing 
Idc464 0 50464 pwl(0 0uA 5ns 14.0680uA) 
Lflux464 50464 0 57.0000pH 
K464 Lg464 Lflux464 1

Cg464 927 0 50.0000fF 
Lg464 927 928 57.0000pH
B464 927 928 10463 jj0 
Cgg464 928 0 50.0000fF
Vmeas464 928 929 0V

*Flux Biasing 
Idc465 0 50465 pwl(0 0uA 5ns 14.0680uA) 
Lflux465 50465 0 57.0000pH 
K465 Lg465 Lflux465 1

Cg465 929 0 50.0000fF 
Lg465 929 930 57.0000pH
B465 929 930 10464 jj0 
Cgg465 930 0 50.0000fF
Vmeas465 930 931 0V

*Flux Biasing 
Idc466 0 50466 pwl(0 0uA 5ns 14.0680uA) 
Lflux466 50466 0 57.0000pH 
K466 Lg466 Lflux466 1

Cg466 931 0 50.0000fF 
Lg466 931 932 57.0000pH
B466 931 932 10465 jj0 
Cgg466 932 0 50.0000fF
Vmeas466 932 933 0V

*Flux Biasing 
Idc467 0 50467 pwl(0 0uA 5ns 14.0680uA) 
Lflux467 50467 0 57.0000pH 
K467 Lg467 Lflux467 1

Cg467 933 0 50.0000fF 
Lg467 933 934 57.0000pH
B467 933 934 10466 jj0 
Cgg467 934 0 50.0000fF
Vmeas467 934 935 0V

*Flux Biasing 
Idc468 0 50468 pwl(0 0uA 5ns 14.0680uA) 
Lflux468 50468 0 57.0000pH 
K468 Lg468 Lflux468 1

Cg468 935 0 50.0000fF 
Lg468 935 936 57.0000pH
B468 935 936 10467 jj0 
Cgg468 936 0 50.0000fF
Vmeas468 936 937 0V

*Flux Biasing 
Idc469 0 50469 pwl(0 0uA 5ns 14.0680uA) 
Lflux469 50469 0 57.0000pH 
K469 Lg469 Lflux469 1

Cg469 937 0 50.0000fF 
Lg469 937 938 57.0000pH
B469 937 938 10468 jj0 
Cgg469 938 0 50.0000fF
Vmeas469 938 939 0V

*Flux Biasing 
Idc470 0 50470 pwl(0 0uA 5ns 14.0680uA) 
Lflux470 50470 0 57.0000pH 
K470 Lg470 Lflux470 1

Cg470 939 0 50.0000fF 
Lg470 939 940 57.0000pH
B470 939 940 10469 jj0 
Cgg470 940 0 50.0000fF
Vmeas470 940 941 0V

*Flux Biasing 
Idc471 0 50471 pwl(0 0uA 5ns 14.0680uA) 
Lflux471 50471 0 57.0000pH 
K471 Lg471 Lflux471 1

Cg471 941 0 50.0000fF 
Lg471 941 942 57.0000pH
B471 941 942 10470 jj0 
Cgg471 942 0 50.0000fF
Vmeas471 942 943 0V

*Flux Biasing 
Idc472 0 50472 pwl(0 0uA 5ns 14.0680uA) 
Lflux472 50472 0 57.0000pH 
K472 Lg472 Lflux472 1

Cg472 943 0 50.0000fF 
Lg472 943 944 57.0000pH
B472 943 944 10471 jj0 
Cgg472 944 0 50.0000fF
Vmeas472 944 945 0V

*Flux Biasing 
Idc473 0 50473 pwl(0 0uA 5ns 14.0680uA) 
Lflux473 50473 0 57.0000pH 
K473 Lg473 Lflux473 1

Cg473 945 0 50.0000fF 
Lg473 945 946 57.0000pH
B473 945 946 10472 jj0 
Cgg473 946 0 50.0000fF
Vmeas473 946 947 0V

*Flux Biasing 
Idc474 0 50474 pwl(0 0uA 5ns 14.0680uA) 
Lflux474 50474 0 57.0000pH 
K474 Lg474 Lflux474 1

Cg474 947 0 50.0000fF 
Lg474 947 948 57.0000pH
B474 947 948 10473 jj0 
Cgg474 948 0 50.0000fF
Vmeas474 948 949 0V

*Flux Biasing 
Idc475 0 50475 pwl(0 0uA 5ns 14.0680uA) 
Lflux475 50475 0 57.0000pH 
K475 Lg475 Lflux475 1

Cg475 949 0 50.0000fF 
Lg475 949 950 57.0000pH
B475 949 950 10474 jj0 
Cgg475 950 0 50.0000fF
Vmeas475 950 951 0V

*Flux Biasing 
Idc476 0 50476 pwl(0 0uA 5ns 14.0680uA) 
Lflux476 50476 0 57.0000pH 
K476 Lg476 Lflux476 1

Cg476 951 0 50.0000fF 
Lg476 951 952 57.0000pH
B476 951 952 10475 jj0 
Cgg476 952 0 50.0000fF
Vmeas476 952 953 0V

*Flux Biasing 
Idc477 0 50477 pwl(0 0uA 5ns 14.0680uA) 
Lflux477 50477 0 57.0000pH 
K477 Lg477 Lflux477 1

Cg477 953 0 50.0000fF 
Lg477 953 954 57.0000pH
B477 953 954 10476 jj0 
Cgg477 954 0 50.0000fF
Vmeas477 954 955 0V

*Flux Biasing 
Idc478 0 50478 pwl(0 0uA 5ns 14.0680uA) 
Lflux478 50478 0 57.0000pH 
K478 Lg478 Lflux478 1

Cg478 955 0 50.0000fF 
Lg478 955 956 57.0000pH
B478 955 956 10477 jj0 
Cgg478 956 0 50.0000fF
Vmeas478 956 957 0V

*Flux Biasing 
Idc479 0 50479 pwl(0 0uA 5ns 14.0680uA) 
Lflux479 50479 0 57.0000pH 
K479 Lg479 Lflux479 1

Cg479 957 0 50.0000fF 
Lg479 957 958 57.0000pH
B479 957 958 10478 jj0 
Cgg479 958 0 50.0000fF
Vmeas479 958 959 0V

*Flux Biasing 
Idc480 0 50480 pwl(0 0uA 5ns 14.0680uA) 
Lflux480 50480 0 57.0000pH 
K480 Lg480 Lflux480 1

Cg480 959 0 50.0000fF 
Lg480 959 960 57.0000pH
B480 959 960 10479 jj0 
Cgg480 960 0 50.0000fF
Vmeas480 960 961 0V

*Flux Biasing 
Idc481 0 50481 pwl(0 0uA 5ns 14.0680uA) 
Lflux481 50481 0 57.0000pH 
K481 Lg481 Lflux481 1

Cg481 961 0 50.0000fF 
Lg481 961 962 57.0000pH
B481 961 962 10480 jj0 
Cgg481 962 0 50.0000fF
Vmeas481 962 963 0V

*Flux Biasing 
Idc482 0 50482 pwl(0 0uA 5ns 14.0680uA) 
Lflux482 50482 0 57.0000pH 
K482 Lg482 Lflux482 1

Cg482 963 0 50.0000fF 
Lg482 963 964 57.0000pH
B482 963 964 10481 jj0 
Cgg482 964 0 50.0000fF
Vmeas482 964 965 0V

*Flux Biasing 
Idc483 0 50483 pwl(0 0uA 5ns 14.0680uA) 
Lflux483 50483 0 57.0000pH 
K483 Lg483 Lflux483 1

Cg483 965 0 50.0000fF 
Lg483 965 966 57.0000pH
B483 965 966 10482 jj0 
Cgg483 966 0 50.0000fF
Vmeas483 966 967 0V

*Flux Biasing 
Idc484 0 50484 pwl(0 0uA 5ns 14.0680uA) 
Lflux484 50484 0 57.0000pH 
K484 Lg484 Lflux484 1

Cg484 967 0 50.0000fF 
Lg484 967 968 57.0000pH
B484 967 968 10483 jj0 
Cgg484 968 0 50.0000fF
Vmeas484 968 969 0V

*Flux Biasing 
Idc485 0 50485 pwl(0 0uA 5ns 14.0680uA) 
Lflux485 50485 0 57.0000pH 
K485 Lg485 Lflux485 1

Cg485 969 0 50.0000fF 
Lg485 969 970 57.0000pH
B485 969 970 10484 jj0 
Cgg485 970 0 50.0000fF
Vmeas485 970 971 0V

*Flux Biasing 
Idc486 0 50486 pwl(0 0uA 5ns 14.0680uA) 
Lflux486 50486 0 57.0000pH 
K486 Lg486 Lflux486 1

Cg486 971 0 50.0000fF 
Lg486 971 972 57.0000pH
B486 971 972 10485 jj0 
Cgg486 972 0 50.0000fF
Vmeas486 972 973 0V

*Flux Biasing 
Idc487 0 50487 pwl(0 0uA 5ns 14.0680uA) 
Lflux487 50487 0 57.0000pH 
K487 Lg487 Lflux487 1

Cg487 973 0 50.0000fF 
Lg487 973 974 57.0000pH
B487 973 974 10486 jj0 
Cgg487 974 0 50.0000fF
Vmeas487 974 975 0V

*Flux Biasing 
Idc488 0 50488 pwl(0 0uA 5ns 14.0680uA) 
Lflux488 50488 0 57.0000pH 
K488 Lg488 Lflux488 1

Cg488 975 0 50.0000fF 
Lg488 975 976 57.0000pH
B488 975 976 10487 jj0 
Cgg488 976 0 50.0000fF
Vmeas488 976 977 0V

*Flux Biasing 
Idc489 0 50489 pwl(0 0uA 5ns 14.0680uA) 
Lflux489 50489 0 57.0000pH 
K489 Lg489 Lflux489 1

Cg489 977 0 50.0000fF 
Lg489 977 978 57.0000pH
B489 977 978 10488 jj0 
Cgg489 978 0 50.0000fF
Vmeas489 978 979 0V

*Flux Biasing 
Idc490 0 50490 pwl(0 0uA 5ns 14.0680uA) 
Lflux490 50490 0 57.0000pH 
K490 Lg490 Lflux490 1

Cg490 979 0 50.0000fF 
Lg490 979 980 57.0000pH
B490 979 980 10489 jj0 
Cgg490 980 0 50.0000fF
Vmeas490 980 981 0V

*Flux Biasing 
Idc491 0 50491 pwl(0 0uA 5ns 14.0680uA) 
Lflux491 50491 0 57.0000pH 
K491 Lg491 Lflux491 1

Cg491 981 0 50.0000fF 
Lg491 981 982 57.0000pH
B491 981 982 10490 jj0 
Cgg491 982 0 50.0000fF
Vmeas491 982 983 0V

*Flux Biasing 
Idc492 0 50492 pwl(0 0uA 5ns 14.0680uA) 
Lflux492 50492 0 57.0000pH 
K492 Lg492 Lflux492 1

Cg492 983 0 50.0000fF 
Lg492 983 984 57.0000pH
B492 983 984 10491 jj0 
Cgg492 984 0 50.0000fF
Vmeas492 984 985 0V

*Flux Biasing 
Idc493 0 50493 pwl(0 0uA 5ns 14.0680uA) 
Lflux493 50493 0 57.0000pH 
K493 Lg493 Lflux493 1

Cg493 985 0 50.0000fF 
Lg493 985 986 57.0000pH
B493 985 986 10492 jj0 
Cgg493 986 0 50.0000fF
Vmeas493 986 987 0V

*Flux Biasing 
Idc494 0 50494 pwl(0 0uA 5ns 14.0680uA) 
Lflux494 50494 0 57.0000pH 
K494 Lg494 Lflux494 1

Cg494 987 0 50.0000fF 
Lg494 987 988 57.0000pH
B494 987 988 10493 jj0 
Cgg494 988 0 50.0000fF
Vmeas494 988 989 0V

*Flux Biasing 
Idc495 0 50495 pwl(0 0uA 5ns 14.0680uA) 
Lflux495 50495 0 57.0000pH 
K495 Lg495 Lflux495 1

Cg495 989 0 50.0000fF 
Lg495 989 990 57.0000pH
B495 989 990 10494 jj0 
Cgg495 990 0 50.0000fF
Vmeas495 990 991 0V

*Flux Biasing 
Idc496 0 50496 pwl(0 0uA 5ns 14.0680uA) 
Lflux496 50496 0 57.0000pH 
K496 Lg496 Lflux496 1

Cg496 991 0 50.0000fF 
Lg496 991 992 57.0000pH
B496 991 992 10495 jj0 
Cgg496 992 0 50.0000fF
Vmeas496 992 993 0V

*Flux Biasing 
Idc497 0 50497 pwl(0 0uA 5ns 14.0680uA) 
Lflux497 50497 0 57.0000pH 
K497 Lg497 Lflux497 1

Cg497 993 0 50.0000fF 
Lg497 993 994 57.0000pH
B497 993 994 10496 jj0 
Cgg497 994 0 50.0000fF
Vmeas497 994 995 0V

*Flux Biasing 
Idc498 0 50498 pwl(0 0uA 5ns 14.0680uA) 
Lflux498 50498 0 57.0000pH 
K498 Lg498 Lflux498 1

Cg498 995 0 50.0000fF 
Lg498 995 996 57.0000pH
B498 995 996 10497 jj0 
Cgg498 996 0 50.0000fF
Vmeas498 996 997 0V

*Flux Biasing 
Idc499 0 50499 pwl(0 0uA 5ns 14.0680uA) 
Lflux499 50499 0 57.0000pH 
K499 Lg499 Lflux499 1

Cg499 997 0 50.0000fF 
Lg499 997 998 57.0000pH
B499 997 998 10498 jj0 
Cgg499 998 0 50.0000fF
Vmeas499 998 999 0V

*Flux Biasing 
Idc500 0 50500 pwl(0 0uA 5ns 14.0680uA) 
Lflux500 50500 0 57.0000pH 
K500 Lg500 Lflux500 1

Cg500 999 0 50.0000fF 
Lg500 999 1000 57.0000pH
B500 999 1000 10499 jj0 
Cgg500 1000 0 50.0000fF
Vmeas500 1000 1001 0V

*Flux Biasing 
Idc501 0 50501 pwl(0 0uA 5ns 14.0680uA) 
Lflux501 50501 0 57.0000pH 
K501 Lg501 Lflux501 1

Cg501 1001 0 50.0000fF 
Lg501 1001 1002 57.0000pH
B501 1001 1002 10500 jj0 
Cgg501 1002 0 50.0000fF
Vmeas501 1002 1003 0V


*Termination Resistor 
Rtermend 1003 0 23.8747Ohm 

.tran 1p 20.0000n 0n uic
.control 
set maxdata = 8e8 
run 

print /printnoheaders time > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/time.txt
print /printnoheaders Vmeas0#branch Vmeas1#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I_initial.txt 

print /printnoheaders v(4) v(6) v(8) v(10) v(12) v(14) v(16) v(18) v(20) v(22) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(1-10).txt 

print /printnoheaders v(24) v(26) v(28) v(30) v(32) v(34) v(36) v(38) v(40) v(42) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(11-20).txt 

print /printnoheaders v(44) v(46) v(48) v(50) v(52) v(54) v(56) v(58) v(60) v(62) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(21-30).txt 

print /printnoheaders v(64) v(66) v(68) v(70) v(72) v(74) v(76) v(78) v(80) v(82) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(31-40).txt 

print /printnoheaders v(84) v(86) v(88) v(90) v(92) v(94) v(96) v(98) v(100) v(102) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(41-50).txt 

print /printnoheaders v(104) v(106) v(108) v(110) v(112) v(114) v(116) v(118) v(120) v(122) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(51-60).txt 

print /printnoheaders v(124) v(126) v(128) v(130) v(132) v(134) v(136) v(138) v(140) v(142) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(61-70).txt 

print /printnoheaders v(144) v(146) v(148) v(150) v(152) v(154) v(156) v(158) v(160) v(162) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(71-80).txt 

print /printnoheaders v(164) v(166) v(168) v(170) v(172) v(174) v(176) v(178) v(180) v(182) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(81-90).txt 

print /printnoheaders v(184) v(186) v(188) v(190) v(192) v(194) v(196) v(198) v(200) v(202) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(91-100).txt 

print /printnoheaders v(204) v(206) v(208) v(210) v(212) v(214) v(216) v(218) v(220) v(222) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(101-110).txt 

print /printnoheaders v(224) v(226) v(228) v(230) v(232) v(234) v(236) v(238) v(240) v(242) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(111-120).txt 

print /printnoheaders v(244) v(246) v(248) v(250) v(252) v(254) v(256) v(258) v(260) v(262) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(121-130).txt 

print /printnoheaders v(264) v(266) v(268) v(270) v(272) v(274) v(276) v(278) v(280) v(282) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(131-140).txt 

print /printnoheaders v(284) v(286) v(288) v(290) v(292) v(294) v(296) v(298) v(300) v(302) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(141-150).txt 

print /printnoheaders v(304) v(306) v(308) v(310) v(312) v(314) v(316) v(318) v(320) v(322) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(151-160).txt 

print /printnoheaders v(324) v(326) v(328) v(330) v(332) v(334) v(336) v(338) v(340) v(342) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(161-170).txt 

print /printnoheaders v(344) v(346) v(348) v(350) v(352) v(354) v(356) v(358) v(360) v(362) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(171-180).txt 

print /printnoheaders v(364) v(366) v(368) v(370) v(372) v(374) v(376) v(378) v(380) v(382) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(181-190).txt 

print /printnoheaders v(384) v(386) v(388) v(390) v(392) v(394) v(396) v(398) v(400) v(402) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(191-200).txt 

print /printnoheaders v(404) v(406) v(408) v(410) v(412) v(414) v(416) v(418) v(420) v(422) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(201-210).txt 

print /printnoheaders v(424) v(426) v(428) v(430) v(432) v(434) v(436) v(438) v(440) v(442) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(211-220).txt 

print /printnoheaders v(444) v(446) v(448) v(450) v(452) v(454) v(456) v(458) v(460) v(462) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(221-230).txt 

print /printnoheaders v(464) v(466) v(468) v(470) v(472) v(474) v(476) v(478) v(480) v(482) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(231-240).txt 

print /printnoheaders v(484) v(486) v(488) v(490) v(492) v(494) v(496) v(498) v(500) v(502) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(241-250).txt 

print /printnoheaders v(504) v(506) v(508) v(510) v(512) v(514) v(516) v(518) v(520) v(522) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(251-260).txt 

print /printnoheaders v(524) v(526) v(528) v(530) v(532) v(534) v(536) v(538) v(540) v(542) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(261-270).txt 

print /printnoheaders v(544) v(546) v(548) v(550) v(552) v(554) v(556) v(558) v(560) v(562) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(271-280).txt 

print /printnoheaders v(564) v(566) v(568) v(570) v(572) v(574) v(576) v(578) v(580) v(582) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(281-290).txt 

print /printnoheaders v(584) v(586) v(588) v(590) v(592) v(594) v(596) v(598) v(600) v(602) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(291-300).txt 

print /printnoheaders v(604) v(606) v(608) v(610) v(612) v(614) v(616) v(618) v(620) v(622) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(301-310).txt 

print /printnoheaders v(624) v(626) v(628) v(630) v(632) v(634) v(636) v(638) v(640) v(642) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(311-320).txt 

print /printnoheaders v(644) v(646) v(648) v(650) v(652) v(654) v(656) v(658) v(660) v(662) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(321-330).txt 

print /printnoheaders v(664) v(666) v(668) v(670) v(672) v(674) v(676) v(678) v(680) v(682) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(331-340).txt 

print /printnoheaders v(684) v(686) v(688) v(690) v(692) v(694) v(696) v(698) v(700) v(702) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(341-350).txt 

print /printnoheaders v(704) v(706) v(708) v(710) v(712) v(714) v(716) v(718) v(720) v(722) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(351-360).txt 

print /printnoheaders v(724) v(726) v(728) v(730) v(732) v(734) v(736) v(738) v(740) v(742) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(361-370).txt 

print /printnoheaders v(744) v(746) v(748) v(750) v(752) v(754) v(756) v(758) v(760) v(762) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(371-380).txt 

print /printnoheaders v(764) v(766) v(768) v(770) v(772) v(774) v(776) v(778) v(780) v(782) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(381-390).txt 

print /printnoheaders v(784) v(786) v(788) v(790) v(792) v(794) v(796) v(798) v(800) v(802) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(391-400).txt 

print /printnoheaders v(804) v(806) v(808) v(810) v(812) v(814) v(816) v(818) v(820) v(822) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(401-410).txt 

print /printnoheaders v(824) v(826) v(828) v(830) v(832) v(834) v(836) v(838) v(840) v(842) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(411-420).txt 

print /printnoheaders v(844) v(846) v(848) v(850) v(852) v(854) v(856) v(858) v(860) v(862) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(421-430).txt 

print /printnoheaders v(864) v(866) v(868) v(870) v(872) v(874) v(876) v(878) v(880) v(882) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(431-440).txt 

print /printnoheaders v(884) v(886) v(888) v(890) v(892) v(894) v(896) v(898) v(900) v(902) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(441-450).txt 

print /printnoheaders v(904) v(906) v(908) v(910) v(912) v(914) v(916) v(918) v(920) v(922) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(451-460).txt 

print /printnoheaders v(924) v(926) v(928) v(930) v(932) v(934) v(936) v(938) v(940) v(942) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(461-470).txt 

print /printnoheaders v(944) v(946) v(948) v(950) v(952) v(954) v(956) v(958) v(960) v(962) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(471-480).txt 

print /printnoheaders v(964) v(966) v(968) v(970) v(972) v(974) v(976) v(978) v(980) v(982) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(481-490).txt 

print /printnoheaders v(984) v(986) v(988) v(990) v(992) v(994) v(996) v(998) v(1000) v(1002) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/V(491-500).txt 

print /printnoheaders v(10001) v(10002) v(10003) v(10004) v(10005) v(10006) v(10007) v(10008) v(10009) v(10010) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10001-10010)-t.txt 

print /printnoheaders v(10011) v(10012) v(10013) v(10014) v(10015) v(10016) v(10017) v(10018) v(10019) v(10020) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10011-10020)-t.txt 

print /printnoheaders v(10021) v(10022) v(10023) v(10024) v(10025) v(10026) v(10027) v(10028) v(10029) v(10030) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10021-10030)-t.txt 

print /printnoheaders v(10031) v(10032) v(10033) v(10034) v(10035) v(10036) v(10037) v(10038) v(10039) v(10040) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10031-10040)-t.txt 

print /printnoheaders v(10041) v(10042) v(10043) v(10044) v(10045) v(10046) v(10047) v(10048) v(10049) v(10050) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10041-10050)-t.txt 

print /printnoheaders v(10051) v(10052) v(10053) v(10054) v(10055) v(10056) v(10057) v(10058) v(10059) v(10060) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10051-10060)-t.txt 

print /printnoheaders v(10061) v(10062) v(10063) v(10064) v(10065) v(10066) v(10067) v(10068) v(10069) v(10070) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10061-10070)-t.txt 

print /printnoheaders v(10071) v(10072) v(10073) v(10074) v(10075) v(10076) v(10077) v(10078) v(10079) v(10080) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10071-10080)-t.txt 

print /printnoheaders v(10081) v(10082) v(10083) v(10084) v(10085) v(10086) v(10087) v(10088) v(10089) v(10090) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10081-10090)-t.txt 

print /printnoheaders v(10091) v(10092) v(10093) v(10094) v(10095) v(10096) v(10097) v(10098) v(10099) v(10100) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10091-10100)-t.txt 

print /printnoheaders v(10101) v(10102) v(10103) v(10104) v(10105) v(10106) v(10107) v(10108) v(10109) v(10110) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10101-10110)-t.txt 

print /printnoheaders v(10111) v(10112) v(10113) v(10114) v(10115) v(10116) v(10117) v(10118) v(10119) v(10120) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10111-10120)-t.txt 

print /printnoheaders v(10121) v(10122) v(10123) v(10124) v(10125) v(10126) v(10127) v(10128) v(10129) v(10130) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10121-10130)-t.txt 

print /printnoheaders v(10131) v(10132) v(10133) v(10134) v(10135) v(10136) v(10137) v(10138) v(10139) v(10140) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10131-10140)-t.txt 

print /printnoheaders v(10141) v(10142) v(10143) v(10144) v(10145) v(10146) v(10147) v(10148) v(10149) v(10150) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10141-10150)-t.txt 

print /printnoheaders v(10151) v(10152) v(10153) v(10154) v(10155) v(10156) v(10157) v(10158) v(10159) v(10160) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10151-10160)-t.txt 

print /printnoheaders v(10161) v(10162) v(10163) v(10164) v(10165) v(10166) v(10167) v(10168) v(10169) v(10170) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10161-10170)-t.txt 

print /printnoheaders v(10171) v(10172) v(10173) v(10174) v(10175) v(10176) v(10177) v(10178) v(10179) v(10180) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10171-10180)-t.txt 

print /printnoheaders v(10181) v(10182) v(10183) v(10184) v(10185) v(10186) v(10187) v(10188) v(10189) v(10190) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10181-10190)-t.txt 

print /printnoheaders v(10191) v(10192) v(10193) v(10194) v(10195) v(10196) v(10197) v(10198) v(10199) v(10200) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10191-10200)-t.txt 

print /printnoheaders v(10201) v(10202) v(10203) v(10204) v(10205) v(10206) v(10207) v(10208) v(10209) v(10210) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10201-10210)-t.txt 

print /printnoheaders v(10211) v(10212) v(10213) v(10214) v(10215) v(10216) v(10217) v(10218) v(10219) v(10220) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10211-10220)-t.txt 

print /printnoheaders v(10221) v(10222) v(10223) v(10224) v(10225) v(10226) v(10227) v(10228) v(10229) v(10230) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10221-10230)-t.txt 

print /printnoheaders v(10231) v(10232) v(10233) v(10234) v(10235) v(10236) v(10237) v(10238) v(10239) v(10240) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10231-10240)-t.txt 

print /printnoheaders v(10241) v(10242) v(10243) v(10244) v(10245) v(10246) v(10247) v(10248) v(10249) v(10250) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10241-10250)-t.txt 

print /printnoheaders v(10251) v(10252) v(10253) v(10254) v(10255) v(10256) v(10257) v(10258) v(10259) v(10260) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10251-10260)-t.txt 

print /printnoheaders v(10261) v(10262) v(10263) v(10264) v(10265) v(10266) v(10267) v(10268) v(10269) v(10270) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10261-10270)-t.txt 

print /printnoheaders v(10271) v(10272) v(10273) v(10274) v(10275) v(10276) v(10277) v(10278) v(10279) v(10280) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10271-10280)-t.txt 

print /printnoheaders v(10281) v(10282) v(10283) v(10284) v(10285) v(10286) v(10287) v(10288) v(10289) v(10290) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10281-10290)-t.txt 

print /printnoheaders v(10291) v(10292) v(10293) v(10294) v(10295) v(10296) v(10297) v(10298) v(10299) v(10300) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10291-10300)-t.txt 

print /printnoheaders v(10301) v(10302) v(10303) v(10304) v(10305) v(10306) v(10307) v(10308) v(10309) v(10310) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10301-10310)-t.txt 

print /printnoheaders v(10311) v(10312) v(10313) v(10314) v(10315) v(10316) v(10317) v(10318) v(10319) v(10320) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10311-10320)-t.txt 

print /printnoheaders v(10321) v(10322) v(10323) v(10324) v(10325) v(10326) v(10327) v(10328) v(10329) v(10330) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10321-10330)-t.txt 

print /printnoheaders v(10331) v(10332) v(10333) v(10334) v(10335) v(10336) v(10337) v(10338) v(10339) v(10340) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10331-10340)-t.txt 

print /printnoheaders v(10341) v(10342) v(10343) v(10344) v(10345) v(10346) v(10347) v(10348) v(10349) v(10350) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10341-10350)-t.txt 

print /printnoheaders v(10351) v(10352) v(10353) v(10354) v(10355) v(10356) v(10357) v(10358) v(10359) v(10360) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10351-10360)-t.txt 

print /printnoheaders v(10361) v(10362) v(10363) v(10364) v(10365) v(10366) v(10367) v(10368) v(10369) v(10370) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10361-10370)-t.txt 

print /printnoheaders v(10371) v(10372) v(10373) v(10374) v(10375) v(10376) v(10377) v(10378) v(10379) v(10380) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10371-10380)-t.txt 

print /printnoheaders v(10381) v(10382) v(10383) v(10384) v(10385) v(10386) v(10387) v(10388) v(10389) v(10390) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10381-10390)-t.txt 

print /printnoheaders v(10391) v(10392) v(10393) v(10394) v(10395) v(10396) v(10397) v(10398) v(10399) v(10400) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10391-10400)-t.txt 

print /printnoheaders v(10401) v(10402) v(10403) v(10404) v(10405) v(10406) v(10407) v(10408) v(10409) v(10410) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10401-10410)-t.txt 

print /printnoheaders v(10411) v(10412) v(10413) v(10414) v(10415) v(10416) v(10417) v(10418) v(10419) v(10420) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10411-10420)-t.txt 

print /printnoheaders v(10421) v(10422) v(10423) v(10424) v(10425) v(10426) v(10427) v(10428) v(10429) v(10430) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10421-10430)-t.txt 

print /printnoheaders v(10431) v(10432) v(10433) v(10434) v(10435) v(10436) v(10437) v(10438) v(10439) v(10440) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10431-10440)-t.txt 

print /printnoheaders v(10441) v(10442) v(10443) v(10444) v(10445) v(10446) v(10447) v(10448) v(10449) v(10450) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10441-10450)-t.txt 

print /printnoheaders v(10451) v(10452) v(10453) v(10454) v(10455) v(10456) v(10457) v(10458) v(10459) v(10460) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10451-10460)-t.txt 

print /printnoheaders v(10461) v(10462) v(10463) v(10464) v(10465) v(10466) v(10467) v(10468) v(10469) v(10470) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10461-10470)-t.txt 

print /printnoheaders v(10471) v(10472) v(10473) v(10474) v(10475) v(10476) v(10477) v(10478) v(10479) v(10480) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10471-10480)-t.txt 

print /printnoheaders v(10481) v(10482) v(10483) v(10484) v(10485) v(10486) v(10487) v(10488) v(10489) v(10490) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10481-10490)-t.txt 

print /printnoheaders v(10491) v(10492) v(10493) v(10494) v(10495) v(10496) v(10497) v(10498) v(10499) v(10500) > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/Phi(10491-10500)-t.txt 

print /printnoheaders Vmeas2#branch Vmeas3#branch Vmeas4#branch Vmeas5#branch Vmeas6#branch Vmeas7#branch Vmeas8#branch Vmeas9#branch Vmeas10#branch Vmeas11#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(1-10).txt 

print /printnoheaders Vmeas12#branch Vmeas13#branch Vmeas14#branch Vmeas15#branch Vmeas16#branch Vmeas17#branch Vmeas18#branch Vmeas19#branch Vmeas20#branch Vmeas21#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(11-20).txt 

print /printnoheaders Vmeas22#branch Vmeas23#branch Vmeas24#branch Vmeas25#branch Vmeas26#branch Vmeas27#branch Vmeas28#branch Vmeas29#branch Vmeas30#branch Vmeas31#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(21-30).txt 

print /printnoheaders Vmeas32#branch Vmeas33#branch Vmeas34#branch Vmeas35#branch Vmeas36#branch Vmeas37#branch Vmeas38#branch Vmeas39#branch Vmeas40#branch Vmeas41#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(31-40).txt 

print /printnoheaders Vmeas42#branch Vmeas43#branch Vmeas44#branch Vmeas45#branch Vmeas46#branch Vmeas47#branch Vmeas48#branch Vmeas49#branch Vmeas50#branch Vmeas51#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(41-50).txt 

print /printnoheaders Vmeas52#branch Vmeas53#branch Vmeas54#branch Vmeas55#branch Vmeas56#branch Vmeas57#branch Vmeas58#branch Vmeas59#branch Vmeas60#branch Vmeas61#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(51-60).txt 

print /printnoheaders Vmeas62#branch Vmeas63#branch Vmeas64#branch Vmeas65#branch Vmeas66#branch Vmeas67#branch Vmeas68#branch Vmeas69#branch Vmeas70#branch Vmeas71#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(61-70).txt 

print /printnoheaders Vmeas72#branch Vmeas73#branch Vmeas74#branch Vmeas75#branch Vmeas76#branch Vmeas77#branch Vmeas78#branch Vmeas79#branch Vmeas80#branch Vmeas81#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(71-80).txt 

print /printnoheaders Vmeas82#branch Vmeas83#branch Vmeas84#branch Vmeas85#branch Vmeas86#branch Vmeas87#branch Vmeas88#branch Vmeas89#branch Vmeas90#branch Vmeas91#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(81-90).txt 

print /printnoheaders Vmeas92#branch Vmeas93#branch Vmeas94#branch Vmeas95#branch Vmeas96#branch Vmeas97#branch Vmeas98#branch Vmeas99#branch Vmeas100#branch Vmeas101#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(91-100).txt 

print /printnoheaders Vmeas102#branch Vmeas103#branch Vmeas104#branch Vmeas105#branch Vmeas106#branch Vmeas107#branch Vmeas108#branch Vmeas109#branch Vmeas110#branch Vmeas111#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(101-110).txt 

print /printnoheaders Vmeas112#branch Vmeas113#branch Vmeas114#branch Vmeas115#branch Vmeas116#branch Vmeas117#branch Vmeas118#branch Vmeas119#branch Vmeas120#branch Vmeas121#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(111-120).txt 

print /printnoheaders Vmeas122#branch Vmeas123#branch Vmeas124#branch Vmeas125#branch Vmeas126#branch Vmeas127#branch Vmeas128#branch Vmeas129#branch Vmeas130#branch Vmeas131#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(121-130).txt 

print /printnoheaders Vmeas132#branch Vmeas133#branch Vmeas134#branch Vmeas135#branch Vmeas136#branch Vmeas137#branch Vmeas138#branch Vmeas139#branch Vmeas140#branch Vmeas141#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(131-140).txt 

print /printnoheaders Vmeas142#branch Vmeas143#branch Vmeas144#branch Vmeas145#branch Vmeas146#branch Vmeas147#branch Vmeas148#branch Vmeas149#branch Vmeas150#branch Vmeas151#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(141-150).txt 

print /printnoheaders Vmeas152#branch Vmeas153#branch Vmeas154#branch Vmeas155#branch Vmeas156#branch Vmeas157#branch Vmeas158#branch Vmeas159#branch Vmeas160#branch Vmeas161#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(151-160).txt 

print /printnoheaders Vmeas162#branch Vmeas163#branch Vmeas164#branch Vmeas165#branch Vmeas166#branch Vmeas167#branch Vmeas168#branch Vmeas169#branch Vmeas170#branch Vmeas171#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(161-170).txt 

print /printnoheaders Vmeas172#branch Vmeas173#branch Vmeas174#branch Vmeas175#branch Vmeas176#branch Vmeas177#branch Vmeas178#branch Vmeas179#branch Vmeas180#branch Vmeas181#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(171-180).txt 

print /printnoheaders Vmeas182#branch Vmeas183#branch Vmeas184#branch Vmeas185#branch Vmeas186#branch Vmeas187#branch Vmeas188#branch Vmeas189#branch Vmeas190#branch Vmeas191#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(181-190).txt 

print /printnoheaders Vmeas192#branch Vmeas193#branch Vmeas194#branch Vmeas195#branch Vmeas196#branch Vmeas197#branch Vmeas198#branch Vmeas199#branch Vmeas200#branch Vmeas201#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(191-200).txt 

print /printnoheaders Vmeas202#branch Vmeas203#branch Vmeas204#branch Vmeas205#branch Vmeas206#branch Vmeas207#branch Vmeas208#branch Vmeas209#branch Vmeas210#branch Vmeas211#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(201-210).txt 

print /printnoheaders Vmeas212#branch Vmeas213#branch Vmeas214#branch Vmeas215#branch Vmeas216#branch Vmeas217#branch Vmeas218#branch Vmeas219#branch Vmeas220#branch Vmeas221#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(211-220).txt 

print /printnoheaders Vmeas222#branch Vmeas223#branch Vmeas224#branch Vmeas225#branch Vmeas226#branch Vmeas227#branch Vmeas228#branch Vmeas229#branch Vmeas230#branch Vmeas231#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(221-230).txt 

print /printnoheaders Vmeas232#branch Vmeas233#branch Vmeas234#branch Vmeas235#branch Vmeas236#branch Vmeas237#branch Vmeas238#branch Vmeas239#branch Vmeas240#branch Vmeas241#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(231-240).txt 

print /printnoheaders Vmeas242#branch Vmeas243#branch Vmeas244#branch Vmeas245#branch Vmeas246#branch Vmeas247#branch Vmeas248#branch Vmeas249#branch Vmeas250#branch Vmeas251#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(241-250).txt 

print /printnoheaders Vmeas252#branch Vmeas253#branch Vmeas254#branch Vmeas255#branch Vmeas256#branch Vmeas257#branch Vmeas258#branch Vmeas259#branch Vmeas260#branch Vmeas261#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(251-260).txt 

print /printnoheaders Vmeas262#branch Vmeas263#branch Vmeas264#branch Vmeas265#branch Vmeas266#branch Vmeas267#branch Vmeas268#branch Vmeas269#branch Vmeas270#branch Vmeas271#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(261-270).txt 

print /printnoheaders Vmeas272#branch Vmeas273#branch Vmeas274#branch Vmeas275#branch Vmeas276#branch Vmeas277#branch Vmeas278#branch Vmeas279#branch Vmeas280#branch Vmeas281#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(271-280).txt 

print /printnoheaders Vmeas282#branch Vmeas283#branch Vmeas284#branch Vmeas285#branch Vmeas286#branch Vmeas287#branch Vmeas288#branch Vmeas289#branch Vmeas290#branch Vmeas291#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(281-290).txt 

print /printnoheaders Vmeas292#branch Vmeas293#branch Vmeas294#branch Vmeas295#branch Vmeas296#branch Vmeas297#branch Vmeas298#branch Vmeas299#branch Vmeas300#branch Vmeas301#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(291-300).txt 

print /printnoheaders Vmeas302#branch Vmeas303#branch Vmeas304#branch Vmeas305#branch Vmeas306#branch Vmeas307#branch Vmeas308#branch Vmeas309#branch Vmeas310#branch Vmeas311#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(301-310).txt 

print /printnoheaders Vmeas312#branch Vmeas313#branch Vmeas314#branch Vmeas315#branch Vmeas316#branch Vmeas317#branch Vmeas318#branch Vmeas319#branch Vmeas320#branch Vmeas321#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(311-320).txt 

print /printnoheaders Vmeas322#branch Vmeas323#branch Vmeas324#branch Vmeas325#branch Vmeas326#branch Vmeas327#branch Vmeas328#branch Vmeas329#branch Vmeas330#branch Vmeas331#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(321-330).txt 

print /printnoheaders Vmeas332#branch Vmeas333#branch Vmeas334#branch Vmeas335#branch Vmeas336#branch Vmeas337#branch Vmeas338#branch Vmeas339#branch Vmeas340#branch Vmeas341#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(331-340).txt 

print /printnoheaders Vmeas342#branch Vmeas343#branch Vmeas344#branch Vmeas345#branch Vmeas346#branch Vmeas347#branch Vmeas348#branch Vmeas349#branch Vmeas350#branch Vmeas351#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(341-350).txt 

print /printnoheaders Vmeas352#branch Vmeas353#branch Vmeas354#branch Vmeas355#branch Vmeas356#branch Vmeas357#branch Vmeas358#branch Vmeas359#branch Vmeas360#branch Vmeas361#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(351-360).txt 

print /printnoheaders Vmeas362#branch Vmeas363#branch Vmeas364#branch Vmeas365#branch Vmeas366#branch Vmeas367#branch Vmeas368#branch Vmeas369#branch Vmeas370#branch Vmeas371#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(361-370).txt 

print /printnoheaders Vmeas372#branch Vmeas373#branch Vmeas374#branch Vmeas375#branch Vmeas376#branch Vmeas377#branch Vmeas378#branch Vmeas379#branch Vmeas380#branch Vmeas381#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(371-380).txt 

print /printnoheaders Vmeas382#branch Vmeas383#branch Vmeas384#branch Vmeas385#branch Vmeas386#branch Vmeas387#branch Vmeas388#branch Vmeas389#branch Vmeas390#branch Vmeas391#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(381-390).txt 

print /printnoheaders Vmeas392#branch Vmeas393#branch Vmeas394#branch Vmeas395#branch Vmeas396#branch Vmeas397#branch Vmeas398#branch Vmeas399#branch Vmeas400#branch Vmeas401#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(391-400).txt 

print /printnoheaders Vmeas402#branch Vmeas403#branch Vmeas404#branch Vmeas405#branch Vmeas406#branch Vmeas407#branch Vmeas408#branch Vmeas409#branch Vmeas410#branch Vmeas411#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(401-410).txt 

print /printnoheaders Vmeas412#branch Vmeas413#branch Vmeas414#branch Vmeas415#branch Vmeas416#branch Vmeas417#branch Vmeas418#branch Vmeas419#branch Vmeas420#branch Vmeas421#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(411-420).txt 

print /printnoheaders Vmeas422#branch Vmeas423#branch Vmeas424#branch Vmeas425#branch Vmeas426#branch Vmeas427#branch Vmeas428#branch Vmeas429#branch Vmeas430#branch Vmeas431#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(421-430).txt 

print /printnoheaders Vmeas432#branch Vmeas433#branch Vmeas434#branch Vmeas435#branch Vmeas436#branch Vmeas437#branch Vmeas438#branch Vmeas439#branch Vmeas440#branch Vmeas441#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(431-440).txt 

print /printnoheaders Vmeas442#branch Vmeas443#branch Vmeas444#branch Vmeas445#branch Vmeas446#branch Vmeas447#branch Vmeas448#branch Vmeas449#branch Vmeas450#branch Vmeas451#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(441-450).txt 

print /printnoheaders Vmeas452#branch Vmeas453#branch Vmeas454#branch Vmeas455#branch Vmeas456#branch Vmeas457#branch Vmeas458#branch Vmeas459#branch Vmeas460#branch Vmeas461#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(451-460).txt 

print /printnoheaders Vmeas462#branch Vmeas463#branch Vmeas464#branch Vmeas465#branch Vmeas466#branch Vmeas467#branch Vmeas468#branch Vmeas469#branch Vmeas470#branch Vmeas471#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(461-470).txt 

print /printnoheaders Vmeas472#branch Vmeas473#branch Vmeas474#branch Vmeas475#branch Vmeas476#branch Vmeas477#branch Vmeas478#branch Vmeas479#branch Vmeas480#branch Vmeas481#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(471-480).txt 

print /printnoheaders Vmeas482#branch Vmeas483#branch Vmeas484#branch Vmeas485#branch Vmeas486#branch Vmeas487#branch Vmeas488#branch Vmeas489#branch Vmeas490#branch Vmeas491#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(481-490).txt 

print /printnoheaders Vmeas492#branch Vmeas493#branch Vmeas494#branch Vmeas495#branch Vmeas496#branch Vmeas497#branch Vmeas498#branch Vmeas499#branch Vmeas500#branch Vmeas501#branch > /home/tom/Documents/WRspice/Outputs/23,Apr2020_16:34/Simulation_sweep/RawData/I(491-500).txt 

.endc
